/*******************************************
****** Wuhan university of technology ******
****** Ruige Lee ******
year: 2019
month: 3
date: 4
hour: 17
minutes: 4
second: 20
********************************************/

module prm_LUTX1_Sp_4_5_4_chk512p1(
	input [3:0] x,
	input [4:0] y,
	input [3:0] z,
	output [511:0] edge_mask_512p1
);

	reg [511:0] edge_mask_reg_512p1;
	assign edge_mask_512p1= edge_mask_reg_512p1;

always @( *) begin
    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011001,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010011000,
13'b101010011001,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001111000,
13'b110001111001,
13'b110010001000,
13'b110010001001,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001001000,
13'b111001001001,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001011000,
13'b111001011001,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001101000,
13'b111001101001,
13'b111001110100,
13'b111001110101,
13'b111001111000,
13'b111001111001,
13'b1000000100110,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1001000100101,
13'b1001000110100,
13'b1001000110101,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100100,
13'b1001001100101,
13'b1001001110100,
13'b1010000100101,
13'b1010000110100,
13'b1010000110101,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001100100,
13'b1010001100101,
13'b1011000100100,
13'b1011000100101,
13'b1011000110100,
13'b1011001000100,
13'b1011001010100,
13'b1100000100100,
13'b1100000110100,
13'b1100001000100: edge_mask_reg_512p1[0] <= 1'b1;
 		default: edge_mask_reg_512p1[0] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001010,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001000,
13'b100111001001,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100110,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110100101,
13'b111110101001,
13'b1000101000100,
13'b1000101000101,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100101,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1011101100100,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1011110010100,
13'b1100101110100,
13'b1100110000100: edge_mask_reg_512p1[1] <= 1'b1;
 		default: edge_mask_reg_512p1[1] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111011001,
13'b110111011010,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101001,
13'b111110101010,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111001001,
13'b111111001010,
13'b1000101000100,
13'b1000101000101,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000101,
13'b1000111000110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000101,
13'b1010101100011,
13'b1010101110011,
13'b1010101110100,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1011101110100,
13'b1011110000100,
13'b1011110010100,
13'b1011110010101,
13'b1011110100100,
13'b1011110100101,
13'b1011110110100,
13'b1100110010100,
13'b1100110100100: edge_mask_reg_512p1[2] <= 1'b1;
 		default: edge_mask_reg_512p1[2] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101011000,
13'b10101011001,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b110100001000,
13'b110100001001,
13'b110100011000,
13'b110100011001,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110011000,
13'b110110011001,
13'b110110101000,
13'b110110101001,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110001000,
13'b111110001001,
13'b111110010101,
13'b111110011000,
13'b111110011001,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010100,
13'b1000110010101,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000100,
13'b1001110000101,
13'b1001110010100,
13'b1001110010101,
13'b1010100100100,
13'b1010100100101,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000100,
13'b1010110000101,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100,
13'b1011110000100,
13'b1100101000100,
13'b1100101010100,
13'b1100101100100: edge_mask_reg_512p1[3] <= 1'b1;
 		default: edge_mask_reg_512p1[3] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001001001,
13'b101000111001,
13'b101001001010,
13'b110000111001,
13'b110000111010: edge_mask_reg_512p1[4] <= 1'b1;
 		default: edge_mask_reg_512p1[4] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010011001,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b11010101000,
13'b11010101001,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b110010111000,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101101000,
13'b111011010101,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000101,
13'b111101000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000101,
13'b1000101000110,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1010011010100,
13'b1010011010101,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1010100110101,
13'b1010101000100,
13'b1010101000101,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1011101000101,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000100,
13'b1100100000101,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100110100,
13'b1100100110101,
13'b1101011110100,
13'b1101100000100,
13'b1101100010100,
13'b1101100100100: edge_mask_reg_512p1[5] <= 1'b1;
 		default: edge_mask_reg_512p1[5] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101001001,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001001,
13'b111111010101,
13'b111111010110,
13'b111111011001,
13'b111111101001,
13'b1000101100100,
13'b1000101100101,
13'b1000101110100,
13'b1000101110101,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100110,
13'b1001101110100,
13'b1001101110101,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100101,
13'b1010110000011,
13'b1010110000100,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1011110010100,
13'b1011110100100,
13'b1011110110100,
13'b1011110110101,
13'b1011111000100,
13'b1011111000101,
13'b1011111010100,
13'b1011111100100,
13'b1100110110100,
13'b1100111000100: edge_mask_reg_512p1[6] <= 1'b1;
 		default: edge_mask_reg_512p1[6] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b101010111001,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b110011001001,
13'b110011001010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110101,
13'b1000100110110,
13'b1001011100101,
13'b1001011100110,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110101,
13'b1001100110110,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100110100,
13'b1011100110101,
13'b1100100000100,
13'b1100100000101,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100110100,
13'b1101100010100,
13'b1101100100100: edge_mask_reg_512p1[7] <= 1'b1;
 		default: edge_mask_reg_512p1[7] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110001100,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b101011111011,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110001100,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001010,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110100111100,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101001100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101011100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101101100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110101111100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110001100,
13'b110110010101,
13'b110110010110,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111010,
13'b110110111011,
13'b111100011010,
13'b111100011011,
13'b111100101010,
13'b111100101011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111010,
13'b111100111011,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101010,
13'b111101101011,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111010,
13'b111101111011,
13'b111110000101,
13'b111110000110,
13'b111110001010,
13'b111110001011,
13'b111110010101,
13'b111110010110,
13'b111110011010,
13'b111110011011,
13'b111110101010,
13'b111110101011,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101001011,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101011010,
13'b1000101011011,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101101010,
13'b1000101101011,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111010,
13'b1000101111011,
13'b1000110000101,
13'b1000110000110,
13'b1001100110110,
13'b1001100110111,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000101,
13'b1001110000110,
13'b1001110010101,
13'b1001110010110,
13'b1010100110110,
13'b1010100110111,
13'b1010101000110,
13'b1010101000111,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101110101,
13'b1010101110110,
13'b1010110000101,
13'b1010110000110,
13'b1010110010101,
13'b1010110010110,
13'b1011101000110,
13'b1011101010101,
13'b1011101010110,
13'b1011101100101,
13'b1011101100110,
13'b1011101110101,
13'b1011101110110,
13'b1011110000101,
13'b1011110000110,
13'b1011110010101,
13'b1011110010110,
13'b1100101010101,
13'b1100101010110,
13'b1100101100101,
13'b1100101100110,
13'b1100101110101,
13'b1100101110110,
13'b1100110000101,
13'b1100110000110: edge_mask_reg_512p1[8] <= 1'b1;
 		default: edge_mask_reg_512p1[8] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110001100,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110001100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011001,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110101111100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110001100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110011100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110101100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111011001,
13'b110111011010,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001001,
13'b111111001010,
13'b111111011001,
13'b111111011010,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010101,
13'b1010101110110,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000100,
13'b1010111000101,
13'b1010111010100,
13'b1010111010101,
13'b1011110000101,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110110100,
13'b1011110110101,
13'b1011111000100,
13'b1011111000101,
13'b1011111010101,
13'b1100110000101,
13'b1100110010101,
13'b1100110100101,
13'b1100110110101,
13'b1100111000101: edge_mask_reg_512p1[9] <= 1'b1;
 		default: edge_mask_reg_512p1[9] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b101001011001,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b110001101001,
13'b110001101010,
13'b110001111001,
13'b110001111010,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b110100001010,
13'b111001111001,
13'b111001111010,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011101001,
13'b111011101010,
13'b1000010000110,
13'b1000010000111,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010111,
13'b1000011011000,
13'b1001010000110,
13'b1001010000111,
13'b1001010010110,
13'b1001010010111,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010111,
13'b1010010000110,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011010110,
13'b1010011010111,
13'b1011010010110,
13'b1011010010111,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010110,
13'b1011011010111,
13'b1100010010110,
13'b1100010010111,
13'b1100010100101,
13'b1100010100110,
13'b1100010100111,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1101010100101,
13'b1101010100110,
13'b1101010110101,
13'b1101010110110,
13'b1101011000101,
13'b1101011000110,
13'b1101011010101,
13'b1101011010110,
13'b1110010100101,
13'b1110010100110,
13'b1110010110101,
13'b1110010110110,
13'b1110011000101,
13'b1110011000110,
13'b1110011010110: edge_mask_reg_512p1[10] <= 1'b1;
 		default: edge_mask_reg_512p1[10] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001111001,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001011001,
13'b111001101001,
13'b1000000100110,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1001000100101,
13'b1001000100110,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1010000100101,
13'b1010000110100,
13'b1010000110101,
13'b1010001000100,
13'b1010001000101,
13'b1011000100100,
13'b1011000100101,
13'b1011000110100,
13'b1011000110101,
13'b1011001000100,
13'b1011001000101,
13'b1100000100100,
13'b1100000100101,
13'b1100000110100,
13'b1100000110101,
13'b1100001000100: edge_mask_reg_512p1[11] <= 1'b1;
 		default: edge_mask_reg_512p1[11] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011010,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010011001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011001,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010001001,
13'b110010001010,
13'b111000101000,
13'b111000101001,
13'b111000110101,
13'b111000110110,
13'b111000111000,
13'b111000111001,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001001000,
13'b111001001001,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001011001,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001101001,
13'b111001110100,
13'b111001110101,
13'b111001111001,
13'b1000000100110,
13'b1000000110100,
13'b1000000110101,
13'b1000001000100,
13'b1000001000101,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1001000100101,
13'b1001000110100,
13'b1001000110101,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010100,
13'b1001001010101,
13'b1001001100101,
13'b1010000110100,
13'b1010000110101,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1011000100100,
13'b1011000110100,
13'b1011001000100,
13'b1011001010100,
13'b1100000100100,
13'b1100000110100,
13'b1100001000100: edge_mask_reg_512p1[12] <= 1'b1;
 		default: edge_mask_reg_512p1[12] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001111000,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001010,
13'b10010001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010101,
13'b110001010110,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001111001,
13'b110001111010,
13'b111000100111,
13'b111000101001,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001101001,
13'b111001101010,
13'b1000000100110,
13'b1000000100111,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010101,
13'b1000001010110,
13'b1001000100101,
13'b1001000100110,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010101,
13'b1010000100101,
13'b1010000100110,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000100,
13'b1011000100100,
13'b1011000100101,
13'b1011000110100,
13'b1011000110101,
13'b1011001000100: edge_mask_reg_512p1[13] <= 1'b1;
 		default: edge_mask_reg_512p1[13] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1110001010,
13'b1110011000,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001000,
13'b100111001001,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000110,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110101001,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000101,
13'b110111000110,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110111001,
13'b111111000101,
13'b111111000110,
13'b111111001001,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101001,
13'b1000111000101,
13'b1000111000110,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100110,
13'b1000111100111,
13'b1001111000101,
13'b1001111000110,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100101,
13'b1001111100110,
13'b1010111000101,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100101,
13'b1010111100110,
13'b1011111100100,
13'b1011111100101,
13'b1100111100100: edge_mask_reg_512p1[14] <= 1'b1;
 		default: edge_mask_reg_512p1[14] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1010001010,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011011,
13'b10001101001,
13'b10001111010,
13'b10010001010,
13'b10010001011,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011011,
13'b10100011100,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111010,
13'b11001111011,
13'b11010001010,
13'b11010001011,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001011,
13'b11100001100,
13'b11100011100,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100010111101,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011001101,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011011101,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010011101,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010101101,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101010111101,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011001101,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011011101,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b110001001010,
13'b110001001011,
13'b110001011010,
13'b110001011011,
13'b110001011100,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001101100,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110001111100,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010001100,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010011100,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010101100,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011001100,
13'b110011011010,
13'b110011011011,
13'b110011011100,
13'b110011101010,
13'b110011101011,
13'b110011101100,
13'b110011111010,
13'b110011111011,
13'b110011111100,
13'b110100001011,
13'b111001001011,
13'b111001011010,
13'b111001011011,
13'b111001101010,
13'b111001101011,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111001111011,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010001100,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010011100,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010101100,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111010111100,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011001100,
13'b111011011010,
13'b111011011011,
13'b111011101010,
13'b111011101011,
13'b1000001111000,
13'b1000001111001,
13'b1000010001000,
13'b1000010001001,
13'b1000010001010,
13'b1000010001011,
13'b1000010011000,
13'b1000010011001,
13'b1000010011010,
13'b1000010011011,
13'b1000010101000,
13'b1000010101001,
13'b1000010101010,
13'b1000010101011,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000010111011,
13'b1000011001001,
13'b1000011001010,
13'b1001001101001,
13'b1001001111000,
13'b1001001111001,
13'b1001010001000,
13'b1001010001001,
13'b1001010011000,
13'b1001010011001,
13'b1001010011010,
13'b1001010101000,
13'b1001010101001,
13'b1001010101010,
13'b1001010111000,
13'b1001010111001,
13'b1001010111010,
13'b1001011001001,
13'b1001011001010,
13'b1010001110111,
13'b1010001111000,
13'b1010001111001,
13'b1010010000111,
13'b1010010001000,
13'b1010010001001,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010101010,
13'b1010010111000,
13'b1010010111001,
13'b1010010111010,
13'b1010011001000,
13'b1010011001001,
13'b1010011001010,
13'b1011001101000,
13'b1011001110111,
13'b1011001111000,
13'b1011001111001,
13'b1011010000111,
13'b1011010001000,
13'b1011010001001,
13'b1011010010111,
13'b1011010011000,
13'b1011010011001,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010110111,
13'b1011010111000,
13'b1011010111001,
13'b1011011001000,
13'b1011011001001,
13'b1100001110111,
13'b1100001111000,
13'b1100010000110,
13'b1100010000111,
13'b1100010001000,
13'b1100010001001,
13'b1100010010110,
13'b1100010010111,
13'b1100010011000,
13'b1100010011001,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010101001,
13'b1100010110111,
13'b1100010111000,
13'b1100010111001,
13'b1100011000111,
13'b1100011001000,
13'b1100011001001,
13'b1101001111000,
13'b1101010000110,
13'b1101010000111,
13'b1101010001000,
13'b1101010010110,
13'b1101010010111,
13'b1101010011000,
13'b1101010011001,
13'b1101010100111,
13'b1101010101000,
13'b1101010101001,
13'b1101010110111,
13'b1101010111000,
13'b1101010111001,
13'b1101011000111,
13'b1101011001000,
13'b1101011001001,
13'b1110010000111,
13'b1110010010111,
13'b1110010011000,
13'b1110010100111,
13'b1110010101000,
13'b1110010101001,
13'b1110010110111,
13'b1110010111000,
13'b1110010111001,
13'b1110011000111,
13'b1110011001000,
13'b1111010010111,
13'b1111010100111,
13'b1111010101000,
13'b1111010110111,
13'b1111010111000,
13'b1111011001000: edge_mask_reg_512p1[15] <= 1'b1;
 		default: edge_mask_reg_512p1[15] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101001,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110001100,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110101,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110001100,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110100,
13'b101110110101,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001001,
13'b101111001010,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110100111100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101001100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101011100,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101101100,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110101111100,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110001100,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110011100,
13'b110110100100,
13'b110110100101,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b111100101010,
13'b111100101011,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111010,
13'b111100111011,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010100,
13'b111110010101,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110100100,
13'b111110100101,
13'b111110101010,
13'b111110101011,
13'b111110111010,
13'b1000100110101,
13'b1000100110110,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101011010,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101101010,
13'b1000101110100,
13'b1000101110101,
13'b1000101111010,
13'b1000110000100,
13'b1000110000101,
13'b1000110010100,
13'b1000110010101,
13'b1000110100100,
13'b1000110100101,
13'b1001101010100,
13'b1001101010101,
13'b1001101100100,
13'b1001101100101,
13'b1001101110100,
13'b1001101110101,
13'b1001110000100,
13'b1001110000101,
13'b1001110010100,
13'b1001110010101,
13'b1001110100100,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010110000100,
13'b1010110000101: edge_mask_reg_512p1[16] <= 1'b1;
 		default: edge_mask_reg_512p1[16] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001010,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011001010,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101001,
13'b11100101010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b101010001000,
13'b101010001001,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b111010101000,
13'b111010101001,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111100001000,
13'b111100001001,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1010010110101,
13'b1010011000100,
13'b1010011000101,
13'b1010011010100,
13'b1010011010101,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1011011000100,
13'b1011011000101,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1100011010100,
13'b1100011100100,
13'b1100011110100,
13'b1101011010100,
13'b1101011100100: edge_mask_reg_512p1[17] <= 1'b1;
 		default: edge_mask_reg_512p1[17] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111010,
13'b10011111011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b101000111001,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1010001100100,
13'b1010001100101,
13'b1010001110100,
13'b1010001110101,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1010010100100,
13'b1010010100101,
13'b1011001100100,
13'b1011001100101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100: edge_mask_reg_512p1[18] <= 1'b1;
 		default: edge_mask_reg_512p1[18] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010101,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100001001,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000100,
13'b110110000101,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110001001,
13'b111110001010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110100,
13'b1000101110101,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100: edge_mask_reg_512p1[19] <= 1'b1;
 		default: edge_mask_reg_512p1[19] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101010,
13'b1101101011,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100101,
13'b11110100110,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100100,
13'b100110100101,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100100,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010011,
13'b110110010100,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110000011,
13'b111110000100,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010011,
13'b111110010100,
13'b111110011001,
13'b111110011010,
13'b111110100011,
13'b111110100100,
13'b111110101001,
13'b111110101010,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1000101110011,
13'b1000101110100,
13'b1000110000011,
13'b1000110000100,
13'b1000110010011,
13'b1000110010100,
13'b1000110100011,
13'b1000110100100,
13'b1001101100011,
13'b1001101100100,
13'b1001101110011,
13'b1001101110100,
13'b1001110000011,
13'b1001110000100,
13'b1001110010011,
13'b1001110010100,
13'b1010101100100,
13'b1010101110100,
13'b1010110000100: edge_mask_reg_512p1[20] <= 1'b1;
 		default: edge_mask_reg_512p1[20] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101010,
13'b11100101011,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101010,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101010,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011001100,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011011100,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011101100,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100001001,
13'b111100001010,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001010,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011010,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011110101,
13'b1100011110110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100101,
13'b1101011100110,
13'b1101011110110,
13'b1110011010110,
13'b1110011100110: edge_mask_reg_512p1[21] <= 1'b1;
 		default: edge_mask_reg_512p1[21] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111010111001,
13'b111010111010,
13'b111011001001,
13'b111011001010,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011001000,
13'b1000011010111,
13'b1000011011000,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1000100100111,
13'b1000100101000,
13'b1001011001000,
13'b1001011010111,
13'b1001011011000,
13'b1001011100111,
13'b1001011101000,
13'b1001011110111,
13'b1001011111000,
13'b1001100000111,
13'b1001100001000,
13'b1001100010111,
13'b1001100011000,
13'b1001100100111,
13'b1010011000111,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1010100100111,
13'b1010100101000,
13'b1011011000111,
13'b1011011010110,
13'b1011011010111,
13'b1011011100110,
13'b1011011100111,
13'b1011011110110,
13'b1011011110111,
13'b1011011111000,
13'b1011100000110,
13'b1011100000111,
13'b1011100001000,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100100111,
13'b1100011000111,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1100100100111,
13'b1101011010111,
13'b1101011100110,
13'b1101011100111,
13'b1101011110110,
13'b1101011110111,
13'b1101100000110,
13'b1101100000111,
13'b1101100010110,
13'b1101100010111,
13'b1110011100110,
13'b1110011110110,
13'b1110100000110,
13'b1110100010110: edge_mask_reg_512p1[22] <= 1'b1;
 		default: edge_mask_reg_512p1[22] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110110,
13'b10010110111,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111010,
13'b11011111011,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010001100,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010011100,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010101100,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011000100,
13'b110011000101,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b111001101001,
13'b111001101010,
13'b111001101011,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011010,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101010,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011010100,
13'b1000011010101,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011010100,
13'b1001011010101,
13'b1010010100101,
13'b1010010110100,
13'b1010010110101,
13'b1010011000100,
13'b1010011000101,
13'b1010011010100,
13'b1010011010101,
13'b1011010110100: edge_mask_reg_512p1[23] <= 1'b1;
 		default: edge_mask_reg_512p1[23] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000110,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100,
13'b1011110000100: edge_mask_reg_512p1[24] <= 1'b1;
 		default: edge_mask_reg_512p1[24] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b111100011001,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111110000110,
13'b111110001001,
13'b111110011001,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1001100100101,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1010100110101,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1011101000100,
13'b1011101000101,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1100101000100,
13'b1100101000101,
13'b1100101010100,
13'b1100101010101,
13'b1100101100100,
13'b1100101100101,
13'b1100101110100,
13'b1101101010100: edge_mask_reg_512p1[25] <= 1'b1;
 		default: edge_mask_reg_512p1[25] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11010011100,
13'b11010101011,
13'b11010101100,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111011,
13'b11101111100,
13'b100010101011,
13'b100010101100,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101000111,
13'b100101001000,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111010,
13'b100101111011,
13'b101010101011,
13'b101010101100,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011101101,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101011111101,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100001101,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100011101,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100101101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111011,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011001010,
13'b110011001011,
13'b110011001100,
13'b110011010110,
13'b110011010111,
13'b110011011010,
13'b110011011011,
13'b110011011100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101010,
13'b110011101011,
13'b110011101100,
13'b110011101101,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110011111100,
13'b110011111101,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100001100,
13'b110100001101,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100011100,
13'b110100011101,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100101100,
13'b110100101101,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110100111100,
13'b110101000110,
13'b110101000111,
13'b110101001010,
13'b110101001011,
13'b110101001100,
13'b110101011010,
13'b110101011011,
13'b110101011100,
13'b110101101010,
13'b110101101011,
13'b111011001010,
13'b111011001011,
13'b111011001100,
13'b111011011010,
13'b111011011011,
13'b111011011100,
13'b111011100110,
13'b111011100111,
13'b111011101010,
13'b111011101011,
13'b111011101100,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111010,
13'b111011111011,
13'b111011111100,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001010,
13'b111100001011,
13'b111100001100,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011010,
13'b111100011011,
13'b111100011100,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101010,
13'b111100101011,
13'b111100101100,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111010,
13'b111100111011,
13'b111100111100,
13'b111101000110,
13'b111101000111,
13'b111101001010,
13'b111101001011,
13'b111101001100,
13'b111101011010,
13'b111101011011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011111011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011010,
13'b1000100011011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000110,
13'b1001100000100,
13'b1001100000101,
13'b1001100010100,
13'b1001100010101,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110101,
13'b1001100110110,
13'b1010100100101,
13'b1010100110101: edge_mask_reg_512p1[26] <= 1'b1;
 		default: edge_mask_reg_512p1[26] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b101001011000,
13'b101001011001,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011111000,
13'b101011111001,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110011,
13'b110001110100,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011111000,
13'b110011111001,
13'b111001101000,
13'b111001110011,
13'b111001110100,
13'b111001111000,
13'b111001111001,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001000,
13'b111010001001,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011000,
13'b111010011001,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101000,
13'b111010101001,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111000,
13'b111010111001,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001000,
13'b111011001001,
13'b111011010011,
13'b111011010100,
13'b111011011000,
13'b1000001110100,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1001010000100,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1011010110100,
13'b1011011000100,
13'b1011011010100,
13'b1011011100100: edge_mask_reg_512p1[27] <= 1'b1;
 		default: edge_mask_reg_512p1[27] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001101001,
13'b101001101010,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b111010001001,
13'b111010001010,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b1000010010110,
13'b1000010010111,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1010010010110,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110101,
13'b1011010100110,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011110101,
13'b1100010110101,
13'b1100011000101,
13'b1100011010101,
13'b1100011100101: edge_mask_reg_512p1[28] <= 1'b1;
 		default: edge_mask_reg_512p1[28] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001001,
13'b100110001010,
13'b101011001001,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010011,
13'b111101010100,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101000100,
13'b1000101010011,
13'b1000101010100,
13'b1001100000011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011: edge_mask_reg_512p1[29] <= 1'b1;
 		default: edge_mask_reg_512p1[29] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001010,
13'b11100001011,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011101001,
13'b111011101010,
13'b1000010000101,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010101010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1001010010100,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011100100,
13'b1010010100100,
13'b1010010100101,
13'b1010010110100,
13'b1010010110101,
13'b1010011000100,
13'b1010011010100: edge_mask_reg_512p1[30] <= 1'b1;
 		default: edge_mask_reg_512p1[30] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111001,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110011001000,
13'b110011001001,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b111011011000,
13'b111011011001,
13'b111011100101,
13'b111011100110,
13'b111011101000,
13'b111011101001,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101011001,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000101,
13'b1000101000110,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000101,
13'b1001101000110,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010101000101,
13'b1010101000110,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100110101,
13'b1100100000100,
13'b1100100010100,
13'b1100100100100: edge_mask_reg_512p1[31] <= 1'b1;
 		default: edge_mask_reg_512p1[31] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110001100,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110001100,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001001,
13'b101111001010,
13'b101111011001,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110101111100,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110001100,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110011100,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110101100,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110110111100,
13'b110111000101,
13'b110111000110,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111011001,
13'b110111011010,
13'b111101011010,
13'b111101011011,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101110011,
13'b111101110100,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110110100,
13'b111110111001,
13'b111110111010,
13'b111110111011,
13'b111111001001,
13'b111111001010,
13'b111111001011,
13'b111111011001,
13'b111111011010,
13'b111111011011,
13'b1000101110011,
13'b1000101110100,
13'b1000110000011,
13'b1000110000100,
13'b1000110010011,
13'b1000110010100,
13'b1000110011010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110011: edge_mask_reg_512p1[32] <= 1'b1;
 		default: edge_mask_reg_512p1[32] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001001,
13'b11110001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100101,
13'b100101100110,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b101011010100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100100,
13'b101101100101,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b110011010100,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100100,
13'b110101100101,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101000,
13'b111011101001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101100100,
13'b111101100101,
13'b111101101001,
13'b1000011100011,
13'b1000011110011,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101100100,
13'b1001100010011,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101010011,
13'b1010100100011,
13'b1010100110011: edge_mask_reg_512p1[33] <= 1'b1;
 		default: edge_mask_reg_512p1[33] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001010,
13'b10011001011,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001011,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b110000110110,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001011100,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001101100,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110001111100,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010001100,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b111000110101,
13'b111000110110,
13'b111000111001,
13'b111000111010,
13'b111000111011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001001001,
13'b111001001010,
13'b111001001011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001011011,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001101001,
13'b111001101010,
13'b111001101011,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111001111011,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010101,
13'b111010011001,
13'b111010011010,
13'b111010101010,
13'b1000000110100,
13'b1000001000100,
13'b1000001000101,
13'b1000001001010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001011010,
13'b1000001100011,
13'b1000001100100,
13'b1000001101010,
13'b1000001110011,
13'b1000001110100,
13'b1000010000011,
13'b1000010000100,
13'b1001001000100,
13'b1001001010100,
13'b1001001100100,
13'b1001001110100,
13'b1001010000100: edge_mask_reg_512p1[34] <= 1'b1;
 		default: edge_mask_reg_512p1[34] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001010,
13'b10011001011,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001011,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b110000110110,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001011100,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001101100,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110001111100,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010001100,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b111000110101,
13'b111000111001,
13'b111000111010,
13'b111001000100,
13'b111001000101,
13'b111001001001,
13'b111001001010,
13'b111001001011,
13'b111001010100,
13'b111001010101,
13'b111001011001,
13'b111001011010,
13'b111001011011,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001101001,
13'b111001101010,
13'b111001101011,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001111001,
13'b111001111010,
13'b111001111011,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010100,
13'b111010010101,
13'b111010011001,
13'b111010011010,
13'b111010101010,
13'b1000001000100,
13'b1000001010011,
13'b1000001010100,
13'b1000001100011,
13'b1000001100100,
13'b1000001101010,
13'b1000001110011,
13'b1000001110100,
13'b1000010000011,
13'b1000010000100,
13'b1001001000011,
13'b1001001000100,
13'b1001001010011,
13'b1001001010100,
13'b1001001100011,
13'b1001001100100,
13'b1001001110011,
13'b1001001110100,
13'b1001010000100: edge_mask_reg_512p1[35] <= 1'b1;
 		default: edge_mask_reg_512p1[35] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111010,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010110,
13'b10010010111,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001011100,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001101100,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110001111100,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010001100,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001001001,
13'b111001001010,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001011011,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001101001,
13'b111001101010,
13'b111001101011,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111001111011,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b1000001010011,
13'b1000001010100,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001101010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001111010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100101,
13'b1001001010100,
13'b1001001100100,
13'b1001001110011,
13'b1001001110100,
13'b1001010000011,
13'b1001010000100,
13'b1001010010011,
13'b1001010010100,
13'b1010001100100,
13'b1010001110100,
13'b1010010000100,
13'b1010010010100: edge_mask_reg_512p1[36] <= 1'b1;
 		default: edge_mask_reg_512p1[36] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000110,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b110000110110,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b111000110101,
13'b111000110110,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b1000000110101,
13'b1000000110110,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1001001000101,
13'b1001001000110,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010010100,
13'b1001010010101,
13'b1010001000110,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1011001010101,
13'b1011001100100,
13'b1011001100101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010101,
13'b1100001100101,
13'b1100001110101,
13'b1100010000101: edge_mask_reg_512p1[37] <= 1'b1;
 		default: edge_mask_reg_512p1[37] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100100,
13'b101110100101,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001001,
13'b101111001010,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100100,
13'b110110100101,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111001001,
13'b110111001010,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110011001,
13'b111110011010,
13'b111110100100,
13'b111110101001,
13'b111110101010,
13'b111110111001,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100011,
13'b1000110100100,
13'b1001101010100,
13'b1001101010101,
13'b1001101100100,
13'b1001101100101,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010011,
13'b1001110010100,
13'b1001110100011,
13'b1001110100100,
13'b1010101100100,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010011,
13'b1010110010100,
13'b1010110100100,
13'b1011101110100,
13'b1011110000100: edge_mask_reg_512p1[38] <= 1'b1;
 		default: edge_mask_reg_512p1[38] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001111000,
13'b1001111001,
13'b10001101000,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001101000,
13'b110001101001,
13'b111000100111,
13'b111000101001,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111001,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001011001,
13'b1000000100110,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000101,
13'b1000001000110,
13'b1001000100101,
13'b1001000100110,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000101,
13'b1010000100101,
13'b1010000110100,
13'b1010000110101,
13'b1010001000101,
13'b1011000100100,
13'b1011000100101,
13'b1011000110100,
13'b1011000110101,
13'b1100000100100,
13'b1100000100101,
13'b1100000110100,
13'b1101000100100: edge_mask_reg_512p1[39] <= 1'b1;
 		default: edge_mask_reg_512p1[39] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110001100,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110001100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001001,
13'b101111001010,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101101100,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110101111100,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110001100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110011100,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b111110101010,
13'b111110111010,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111010,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110001010,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1001101010100,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100100,
13'b1010110100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1011110010101,
13'b1011110100101,
13'b1100110010101: edge_mask_reg_512p1[40] <= 1'b1;
 		default: edge_mask_reg_512p1[40] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001010,
13'b10100001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b110001011010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111010,
13'b111001101001,
13'b111001101010,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1100010010100,
13'b1100010010101,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100011000101,
13'b1101010100101,
13'b1101010110101,
13'b1101010110110,
13'b1101011000101: edge_mask_reg_512p1[41] <= 1'b1;
 		default: edge_mask_reg_512p1[41] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001010,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b110100010100,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b111100010100,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101111001,
13'b111110000100,
13'b111110001001,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110011,
13'b1000101110100,
13'b1001100110011,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1001101110011,
13'b1001101110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100,
13'b1010101110011,
13'b1010101110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[42] <= 1'b1;
 		default: edge_mask_reg_512p1[42] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b101001101000,
13'b101001101001,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100001000,
13'b101100001001,
13'b110001111000,
13'b110001111001,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110011,
13'b110011111000,
13'b110011111001,
13'b111001111000,
13'b111001111001,
13'b111010000100,
13'b111010000101,
13'b111010001000,
13'b111010001001,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011000,
13'b111010011001,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101000,
13'b111010101001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111000,
13'b111010111001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001000,
13'b111011001001,
13'b111011010011,
13'b111011010100,
13'b111011011000,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011101000,
13'b111011101001,
13'b1000010000100,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100,
13'b1011011010100: edge_mask_reg_512p1[43] <= 1'b1;
 		default: edge_mask_reg_512p1[43] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001010,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110001100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110001100,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110110101,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001001,
13'b101111001010,
13'b101111011001,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101101100,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110101111100,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110001100,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110011100,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110101100,
13'b110110110101,
13'b110110110110,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111011001,
13'b110111011010,
13'b111101001010,
13'b111101001011,
13'b111101011010,
13'b111101011011,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110111001,
13'b111110111010,
13'b111110111011,
13'b111111001001,
13'b111111001010,
13'b111111001011,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110001010,
13'b1000110001011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110011010,
13'b1000110011011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110101010,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000100,
13'b1001101110110,
13'b1001101110111,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110100,
13'b1001110110101,
13'b1001111000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110100,
13'b1010110110101,
13'b1011110000101,
13'b1011110010100,
13'b1011110010101,
13'b1011110100101,
13'b1011110110101: edge_mask_reg_512p1[44] <= 1'b1;
 		default: edge_mask_reg_512p1[44] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b100011101000,
13'b100011101001,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b101011101000,
13'b101011101001,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b110011111000,
13'b110011111001,
13'b110100000011,
13'b110100000100,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010011,
13'b110100010100,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b111100001000,
13'b111100001001,
13'b111100010011,
13'b111100010100,
13'b111100011000,
13'b111100011001,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011000,
13'b111101011001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101000,
13'b111101101001,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101111001,
13'b111110000011,
13'b111110001001,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000011,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101110011,
13'b1001101110100,
13'b1001110000011,
13'b1010101000011,
13'b1010101010011,
13'b1010101100011,
13'b1010101110011,
13'b1010101110100: edge_mask_reg_512p1[45] <= 1'b1;
 		default: edge_mask_reg_512p1[45] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p1[46] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100101,
13'b11001100110,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001010,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001001,
13'b100100001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100100,
13'b101001100101,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b110001011001,
13'b110001011010,
13'b110001100100,
13'b110001100101,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001100100,
13'b111001101001,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001111001,
13'b111001111010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b1000001110011,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010100,
13'b1000011010101,
13'b1001010000011,
13'b1001010000100,
13'b1001010010011,
13'b1001010010100,
13'b1001010100011,
13'b1001010100100,
13'b1001010110011,
13'b1001010110100,
13'b1001011000011,
13'b1001011000100,
13'b1010010000011,
13'b1010010010011,
13'b1010010010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100: edge_mask_reg_512p1[47] <= 1'b1;
 		default: edge_mask_reg_512p1[47] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001001,
13'b101111001010,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001000,
13'b111101001001,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110101001,
13'b1000100010100,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010100,
13'b1010110010101,
13'b1011101100100,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110010100,
13'b1100101110100,
13'b1100110000100: edge_mask_reg_512p1[48] <= 1'b1;
 		default: edge_mask_reg_512p1[48] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010111001,
13'b1011001000,
13'b1011001001,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100101001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b100001100111,
13'b100001101000,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b101001100111,
13'b101001101000,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b110001110111,
13'b110001111000,
13'b110010000111,
13'b110010001000,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b1000010010101,
13'b1000010010110,
13'b1000010100101,
13'b1000010100110,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110101,
13'b1001010110110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100101,
13'b1001011100110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100101,
13'b1010011100110,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011100101,
13'b1011011100110,
13'b1100010010100,
13'b1100010010101,
13'b1100010100100,
13'b1100010100101,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1101010100100,
13'b1101010100101,
13'b1101010110100,
13'b1101010110101,
13'b1101011000100,
13'b1101011000101,
13'b1101011010100,
13'b1101011010101,
13'b1101011100100,
13'b1101011100101,
13'b1110010110100,
13'b1110011000100,
13'b1110011000101,
13'b1110011010100,
13'b1110011010101,
13'b1110011100100: edge_mask_reg_512p1[49] <= 1'b1;
 		default: edge_mask_reg_512p1[49] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001010,
13'b1001111001,
13'b1010001010,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b10001101000,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b110001001001,
13'b110001001010,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b111001011001,
13'b111001011010,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011001001,
13'b111011001010,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1001001110101,
13'b1001001110110,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1010001110101,
13'b1010001110110,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110100,
13'b1010010110101,
13'b1011001110110,
13'b1011010000101,
13'b1011010000110,
13'b1011010000111,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101,
13'b1100010010110,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010110100,
13'b1100010110101,
13'b1100011000101,
13'b1101010010101,
13'b1101010100101,
13'b1101010100110,
13'b1101010110101: edge_mask_reg_512p1[50] <= 1'b1;
 		default: edge_mask_reg_512p1[50] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111010,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111011,
13'b10001111010,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011010,
13'b100011011011,
13'b100011101010,
13'b100011101011,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011010,
13'b101011011011,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001011100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001101100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110001111100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010001100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010011100,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010101100,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011010,
13'b110011011011,
13'b111000111010,
13'b111000111011,
13'b111001000110,
13'b111001001010,
13'b111001001011,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011010,
13'b111001011011,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101010,
13'b111001101011,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111010,
13'b111001111011,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100110,
13'b111010101010,
13'b111010101011,
13'b111010111010,
13'b111010111011,
13'b111011001010,
13'b111011001011,
13'b1000001000110,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001101010,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000001111010,
13'b1000001111011,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010001010,
13'b1000010001011,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010011011,
13'b1000010100110,
13'b1000010100111,
13'b1001001000110,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1010001010110,
13'b1010001010111,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010100101,
13'b1010010100110,
13'b1010010110101,
13'b1010010110110,
13'b1011001100101,
13'b1011001100110,
13'b1011001110101,
13'b1011001110110,
13'b1011010000101,
13'b1011010000110,
13'b1011010000111,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010100101,
13'b1011010100110,
13'b1011010110101,
13'b1011010110110,
13'b1100001110101,
13'b1100010000101,
13'b1100010000110,
13'b1100010010101,
13'b1100010010110,
13'b1100010100101,
13'b1100010100110,
13'b1100010110110: edge_mask_reg_512p1[51] <= 1'b1;
 		default: edge_mask_reg_512p1[51] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p1[52] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111010,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b110100010101,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101001,
13'b110110101010,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b111110011010,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1010100100100,
13'b1010100110100,
13'b1010100110101,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1010110000100,
13'b1011100110100,
13'b1011101000100,
13'b1011101000101,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1100101100101,
13'b1100101110101: edge_mask_reg_512p1[53] <= 1'b1;
 		default: edge_mask_reg_512p1[53] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001010,
13'b11100001011,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001010,
13'b110001101001,
13'b110001101010,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011101001,
13'b111011101010,
13'b1000010000101,
13'b1000010000110,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1001010000101,
13'b1001010000110,
13'b1001010010101,
13'b1001010010110,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1010010010101,
13'b1010010010110,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010101,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011010101,
13'b1100010100100,
13'b1100010100101,
13'b1100010110100,
13'b1100010110101,
13'b1100011000101,
13'b1100011010101,
13'b1101010110101,
13'b1101011000101: edge_mask_reg_512p1[54] <= 1'b1;
 		default: edge_mask_reg_512p1[54] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10110001001,
13'b10110001010,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000101,
13'b101111000110,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101011001,
13'b110101011010,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000101,
13'b110111000110,
13'b110111001001,
13'b110111001010,
13'b110111011001,
13'b110111011010,
13'b111101001001,
13'b111101001010,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110110100,
13'b111110110101,
13'b111110111001,
13'b111110111010,
13'b111111000100,
13'b111111000101,
13'b111111001001,
13'b111111001010,
13'b1000101010101,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110100,
13'b1000110110101,
13'b1001101100011,
13'b1001101100100,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110100011,
13'b1001110100100,
13'b1001110110100,
13'b1010101100100,
13'b1010101110100,
13'b1010110000100,
13'b1010110010100,
13'b1010110100100,
13'b1011101110100,
13'b1011110000100: edge_mask_reg_512p1[55] <= 1'b1;
 		default: edge_mask_reg_512p1[55] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011111001,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101011000,
13'b100101011001,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101011000,
13'b101101011001,
13'b110011001000,
13'b110011001001,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101011000,
13'b110101011001,
13'b111011011000,
13'b111011100101,
13'b111011100110,
13'b111011101000,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110101,
13'b111100110110,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1010100110101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1100011110100,
13'b1100100000100,
13'b1100100010100: edge_mask_reg_512p1[56] <= 1'b1;
 		default: edge_mask_reg_512p1[56] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101011,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010011100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010101100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011001100,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011011100,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011101100,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011010,
13'b110100011011,
13'b111001101001,
13'b111001101010,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011111010,
13'b111011111011,
13'b111100001010,
13'b1000010000101,
13'b1000010000110,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001010,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011010,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1001010000101,
13'b1001010000110,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1011010010110,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1100010100101,
13'b1100010100110,
13'b1100010110101,
13'b1100010110110,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011100101,
13'b1100011100110,
13'b1101010100101,
13'b1101010110101,
13'b1101010110110,
13'b1101011000101,
13'b1101011000110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100110: edge_mask_reg_512p1[57] <= 1'b1;
 		default: edge_mask_reg_512p1[57] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010101,
13'b101110010110,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101001,
13'b111110101010,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000110010101,
13'b1000110010110,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100110,
13'b1001110010101,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100101,
13'b1001111100110,
13'b1010110100100,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111010100,
13'b1010111010101,
13'b1011110110100,
13'b1011111000100,
13'b1011111010100: edge_mask_reg_512p1[58] <= 1'b1;
 		default: edge_mask_reg_512p1[58] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001011001,
13'b11001011010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b111000100111,
13'b111000101001,
13'b111000110101,
13'b111000111001,
13'b1000000100110,
13'b1000000110101,
13'b1001000100101,
13'b1001000100110: edge_mask_reg_512p1[59] <= 1'b1;
 		default: edge_mask_reg_512p1[59] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001010,
13'b10010001011,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111010,
13'b11011111011,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111010,
13'b100011111011,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111010,
13'b101011111011,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101010,
13'b110011101011,
13'b110011111011,
13'b111001001010,
13'b111001001011,
13'b111001011010,
13'b111001011011,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001101011,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111001111011,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011001010,
13'b111011001011,
13'b111011011010,
13'b111011011011,
13'b1000001100111,
13'b1000001101000,
13'b1000001101001,
13'b1000001110111,
13'b1000001111000,
13'b1000001111001,
13'b1000001111010,
13'b1000010000111,
13'b1000010001000,
13'b1000010001001,
13'b1000010001010,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010011010,
13'b1000010011011,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010101010,
13'b1000010101011,
13'b1000010111000,
13'b1000010111001,
13'b1000011001000,
13'b1001001100111,
13'b1001001101000,
13'b1001001110111,
13'b1001001111000,
13'b1001010000111,
13'b1001010001000,
13'b1001010001001,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1010001100111,
13'b1010001101000,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110111,
13'b1010010111000,
13'b1010011001000,
13'b1011001100111,
13'b1011001101000,
13'b1011001110110,
13'b1011001110111,
13'b1011001111000,
13'b1011010000110,
13'b1011010000111,
13'b1011010001000,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1100001100111,
13'b1100001110110,
13'b1100001110111,
13'b1100001111000,
13'b1100010000110,
13'b1100010000111,
13'b1100010001000,
13'b1100010010110,
13'b1100010010111,
13'b1100010011000,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1101001110110,
13'b1101010000110,
13'b1101010000111,
13'b1101010010110,
13'b1101010010111,
13'b1101010100110,
13'b1101010100111,
13'b1101010101000,
13'b1101010110110,
13'b1101010110111,
13'b1110010000110,
13'b1110010010110,
13'b1110010100110,
13'b1110010100111,
13'b1110010110110: edge_mask_reg_512p1[60] <= 1'b1;
 		default: edge_mask_reg_512p1[60] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101101001,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110101001,
13'b111110101010,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b1000110110110,
13'b1000110110111,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110110110,
13'b1001110110111,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1011111000101,
13'b1011111000110,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1011111110111,
13'b1100111000101,
13'b1100111000110,
13'b1100111010101,
13'b1100111010110,
13'b1100111100101,
13'b1100111100110,
13'b1100111110101,
13'b1100111110110,
13'b1101111000101,
13'b1101111000110,
13'b1101111010101,
13'b1101111010110,
13'b1101111100101,
13'b1101111100110,
13'b1101111110101: edge_mask_reg_512p1[61] <= 1'b1;
 		default: edge_mask_reg_512p1[61] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001010,
13'b10100001011,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001011001,
13'b111001011010,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1010001110110,
13'b1010010000101,
13'b1010010000110,
13'b1010010010101,
13'b1010010010110,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110101,
13'b1010010110110,
13'b1010011000101,
13'b1010011000110,
13'b1011010010101,
13'b1011010010110,
13'b1011010100101,
13'b1011010100110,
13'b1011010110101,
13'b1011010110110,
13'b1011011000101,
13'b1011011000110,
13'b1011011010101,
13'b1100010100101,
13'b1100010110101,
13'b1100011000101,
13'b1100011010101,
13'b1101010110101,
13'b1101011000101: edge_mask_reg_512p1[62] <= 1'b1;
 		default: edge_mask_reg_512p1[62] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001010,
13'b11011001011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001010,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001001001,
13'b111001001010,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010101,
13'b1001001000101,
13'b1001001000110,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010100,
13'b1001010010101,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1100001100100,
13'b1100001100101,
13'b1100001110100,
13'b1100001110101,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101,
13'b1101001110100: edge_mask_reg_512p1[63] <= 1'b1;
 		default: edge_mask_reg_512p1[63] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011010,
13'b11100011011,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b101001101010,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b111010001001,
13'b111010001010,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b1000010010110,
13'b1000010010111,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100110,
13'b1000011100111,
13'b1001010010110,
13'b1001010010111,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100110,
13'b1001011100111,
13'b1010010010110,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100110,
13'b1011010100110,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1100010110101,
13'b1100010110110,
13'b1100011000101,
13'b1100011000110,
13'b1100011010101,
13'b1100011010110,
13'b1100011100101,
13'b1101011000101,
13'b1101011010101: edge_mask_reg_512p1[64] <= 1'b1;
 		default: edge_mask_reg_512p1[64] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110000111,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110001100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110001100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101101010,
13'b110101101011,
13'b110101101100,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110101111100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110001100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110011100,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110101100,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110110111100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011001,
13'b110111011010,
13'b111101111010,
13'b111101111011,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001010,
13'b111110001011,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011010,
13'b111110011011,
13'b111110011100,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101010,
13'b111110101011,
13'b111110101100,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111010,
13'b111110111011,
13'b111110111100,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001010,
13'b111111001011,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011010,
13'b111111011011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110101010,
13'b1000110101011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000110111010,
13'b1000110111011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111001010,
13'b1000111001011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1001110010100,
13'b1001110010101,
13'b1001110100100,
13'b1001110100101,
13'b1001110110100,
13'b1001110110101,
13'b1001111000100,
13'b1001111000101,
13'b1001111010100,
13'b1001111010101,
13'b1010110100101,
13'b1010110110101,
13'b1010111000101: edge_mask_reg_512p1[65] <= 1'b1;
 		default: edge_mask_reg_512p1[65] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110100011001,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b111110101010,
13'b1000101000100,
13'b1000101000101,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1001101000101,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1100101100100,
13'b1100101100101,
13'b1100101110100,
13'b1100101110101,
13'b1100110000100,
13'b1100110000101: edge_mask_reg_512p1[66] <= 1'b1;
 		default: edge_mask_reg_512p1[66] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101010,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111000,
13'b110110111001,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101001000,
13'b111101001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010100,
13'b111110010101,
13'b111110011001,
13'b111110101001,
13'b1000101000100,
13'b1000101000101,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010011,
13'b1001110010100,
13'b1001110100011,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010011,
13'b1010110010100,
13'b1010110100011,
13'b1011101100100,
13'b1011101110100,
13'b1011110000100,
13'b1011110010100,
13'b1100101100100,
13'b1100101110100: edge_mask_reg_512p1[67] <= 1'b1;
 		default: edge_mask_reg_512p1[67] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110100001010,
13'b111001101001,
13'b111001101010,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011101001,
13'b111011101010,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1001010000101,
13'b1001010000110,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010100,
13'b1001011010101,
13'b1001011100100,
13'b1001011100101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000100,
13'b1010011000101,
13'b1010011010100,
13'b1010011010101,
13'b1010011100100,
13'b1010011100101,
13'b1011010100101,
13'b1011010110100,
13'b1011010110101,
13'b1011011000100,
13'b1011011000101,
13'b1011011010100,
13'b1011011010101,
13'b1011011100101: edge_mask_reg_512p1[68] <= 1'b1;
 		default: edge_mask_reg_512p1[68] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101101011001,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101111001,
13'b111101111010,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110000110,
13'b1001110000111,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100110,
13'b1001111100111,
13'b1010110000110,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1011110000110,
13'b1011110010101,
13'b1011110010110,
13'b1011110100101,
13'b1011110100110,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1100110010101,
13'b1100110100101,
13'b1100110100110,
13'b1100110110101,
13'b1100110110110,
13'b1100111000101,
13'b1100111000110,
13'b1100111010101,
13'b1100111010110,
13'b1100111100101,
13'b1100111100110,
13'b1101110010101,
13'b1101110100101,
13'b1101110110101,
13'b1101111000101,
13'b1101111010101,
13'b1101111100101: edge_mask_reg_512p1[69] <= 1'b1;
 		default: edge_mask_reg_512p1[69] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110001100,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110001100,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001010,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101011100,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101101100,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110101111100,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110001100,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110011100,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111001010,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b1000101000110,
13'b1000101000111,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000101111010,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110010111,
13'b1000110011000,
13'b1001101000110,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010111,
13'b1010101010110,
13'b1010101010111,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110010110,
13'b1010110010111,
13'b1011101010110,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1011101110101,
13'b1011101110110,
13'b1011101110111,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110010101,
13'b1011110010110,
13'b1100101100101,
13'b1100101100110,
13'b1100101110101,
13'b1100101110110,
13'b1100110000101,
13'b1100110000110,
13'b1100110010101,
13'b1100110010110,
13'b1101101110101,
13'b1101101110110,
13'b1101110000101,
13'b1101110000110: edge_mask_reg_512p1[70] <= 1'b1;
 		default: edge_mask_reg_512p1[70] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b10001100110,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111001,
13'b11010111010,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111001,
13'b100010111010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111001,
13'b101010111010,
13'b110000110110,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b111000101001,
13'b111000110101,
13'b111000110110,
13'b111000111001,
13'b111000111010,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010011001,
13'b111010011010,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000010000100,
13'b1000010000101,
13'b1001000110101,
13'b1001001000100,
13'b1001001000101,
13'b1001001010100,
13'b1001001010101,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001010000011,
13'b1001010000100,
13'b1010001000100,
13'b1010001010100,
13'b1010001010101,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001110011,
13'b1010001110100,
13'b1010010000011,
13'b1010010000100,
13'b1010010010100,
13'b1011001010100,
13'b1011001100100,
13'b1011001100101,
13'b1011001110100,
13'b1011010000100: edge_mask_reg_512p1[71] <= 1'b1;
 		default: edge_mask_reg_512p1[71] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b10100011011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001010,
13'b110100001011,
13'b111001011010,
13'b111001011011,
13'b111001101010,
13'b111001101011,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111001111011,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101010,
13'b111011101011,
13'b111011111010,
13'b1000001111000,
13'b1000001111001,
13'b1000010000111,
13'b1000010001000,
13'b1000010001001,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010011010,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010101010,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011001000,
13'b1000011001001,
13'b1000011011000,
13'b1001001111000,
13'b1001010000111,
13'b1001010001000,
13'b1001010001001,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011001000,
13'b1001011001001,
13'b1001011011000,
13'b1010001110111,
13'b1010001111000,
13'b1010010000111,
13'b1010010001000,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010111,
13'b1010011011000,
13'b1011001110111,
13'b1011001111000,
13'b1011010000111,
13'b1011010001000,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110111,
13'b1011010111000,
13'b1011011000111,
13'b1011011001000,
13'b1011011010111,
13'b1011011011000,
13'b1100001110111,
13'b1100001111000,
13'b1100010000111,
13'b1100010001000,
13'b1100010010110,
13'b1100010010111,
13'b1100010011000,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010111,
13'b1100011011000,
13'b1101010000111,
13'b1101010001000,
13'b1101010010110,
13'b1101010010111,
13'b1101010011000,
13'b1101010100110,
13'b1101010100111,
13'b1101010101000,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1110010010110,
13'b1110010010111,
13'b1110010100110,
13'b1110010100111,
13'b1110010110110,
13'b1110010110111,
13'b1110011000110,
13'b1110011000111,
13'b1111010110110,
13'b1111010110111,
13'b1111011000110: edge_mask_reg_512p1[72] <= 1'b1;
 		default: edge_mask_reg_512p1[72] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001001,
13'b101011001010,
13'b110000111001,
13'b110000111010,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b111000111001,
13'b111000111010,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001001011,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001011011,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001101011,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111001111011,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b1000001000111,
13'b1000001001000,
13'b1000001001001,
13'b1000001010111,
13'b1000001011000,
13'b1000001011001,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001101001,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000001111001,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1001001000111,
13'b1001001001000,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1010001000110,
13'b1010001000111,
13'b1010001001000,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1010001100110,
13'b1010001100111,
13'b1010001101000,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010010110,
13'b1010010010111,
13'b1011001000110,
13'b1011001000111,
13'b1011001001000,
13'b1011001010110,
13'b1011001010111,
13'b1011001011000,
13'b1011001100110,
13'b1011001100111,
13'b1011001101000,
13'b1011001110110,
13'b1011001110111,
13'b1011001111000,
13'b1011010000110,
13'b1011010000111,
13'b1011010001000,
13'b1011010010110,
13'b1011010010111,
13'b1100001000111,
13'b1100001010110,
13'b1100001010111,
13'b1100001011000,
13'b1100001100110,
13'b1100001100111,
13'b1100001101000,
13'b1100001110110,
13'b1100001110111,
13'b1100001111000,
13'b1100010000110,
13'b1100010000111,
13'b1100010010110,
13'b1100010010111,
13'b1101001000111,
13'b1101001010111,
13'b1101001011000,
13'b1101001100110,
13'b1101001100111,
13'b1101001101000,
13'b1101001110110,
13'b1101001110111,
13'b1101010000110,
13'b1101010000111,
13'b1101010010110,
13'b1101010010111,
13'b1101010100110,
13'b1110001010111,
13'b1110001100110,
13'b1110001100111,
13'b1110001110110,
13'b1110001110111,
13'b1110010000110,
13'b1110010000111,
13'b1110010010110,
13'b1110010010111,
13'b1110010100110,
13'b1111001100110,
13'b1111001100111,
13'b1111001110110,
13'b1111001110111,
13'b1111010000110,
13'b1111010000111,
13'b1111010010110,
13'b1111010010111,
13'b1111010100110: edge_mask_reg_512p1[73] <= 1'b1;
 		default: edge_mask_reg_512p1[73] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100011010,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000101,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100100,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101000100,
13'b1000101010011,
13'b1001100000011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1010100010011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011: edge_mask_reg_512p1[74] <= 1'b1;
 		default: edge_mask_reg_512p1[74] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001010,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001011,
13'b10001101001,
13'b10001111010,
13'b10010001010,
13'b10010001011,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111011,
13'b10011111100,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101010,
13'b11011101011,
13'b11011111011,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101010,
13'b100011101011,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101010,
13'b101011101011,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001101100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110001111100,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010001100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010011100,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010101100,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011010,
13'b110011011011,
13'b110011101010,
13'b110011101011,
13'b111001001010,
13'b111001001011,
13'b111001011010,
13'b111001011011,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101010,
13'b111001101011,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111010,
13'b111001111011,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010111010,
13'b111010111011,
13'b111011001010,
13'b111011001011,
13'b111011011010,
13'b111011011011,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010011010,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010101010,
13'b1000010110110,
13'b1001001100110,
13'b1001001100111,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1010001100110,
13'b1010001100111,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110110,
13'b1010010110111,
13'b1011001110110,
13'b1011001110111,
13'b1011010000101,
13'b1011010000110,
13'b1011010000111,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010110101,
13'b1011010110110,
13'b1011011000110,
13'b1100010000101,
13'b1100010000110,
13'b1100010010101,
13'b1100010010110,
13'b1100010100101,
13'b1100010100110,
13'b1100010100111,
13'b1100010110101,
13'b1100010110110,
13'b1100011000110,
13'b1101010010110,
13'b1101010100110,
13'b1101010110110: edge_mask_reg_512p1[75] <= 1'b1;
 		default: edge_mask_reg_512p1[75] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b10100011011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b110001011010,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010011100,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010101100,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011001100,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001010,
13'b111001101001,
13'b111001101010,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011111010,
13'b1000010000101,
13'b1000010000110,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101010,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111010,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011001010,
13'b1000011010100,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010100,
13'b1001011010101,
13'b1001011100100,
13'b1001011100101,
13'b1010010100101,
13'b1010010110100,
13'b1010010110101,
13'b1010011000100,
13'b1010011000101,
13'b1010011010100,
13'b1010011010101,
13'b1010011100100,
13'b1010011100101,
13'b1011010110100: edge_mask_reg_512p1[76] <= 1'b1;
 		default: edge_mask_reg_512p1[76] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b1110001010,
13'b10100001011,
13'b10100001100,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11100011011,
13'b11100011100,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110001100,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101101101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101101111101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110001100,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001001,
13'b101111001010,
13'b110100101011,
13'b110100111010,
13'b110100111011,
13'b110100111100,
13'b110101001010,
13'b110101001011,
13'b110101001100,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011010,
13'b110101011011,
13'b110101011100,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101101100,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110101111100,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110001100,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110011100,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110101100,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110110111100,
13'b110111001010,
13'b110111001011,
13'b110111011010,
13'b111100111011,
13'b111101001010,
13'b111101001011,
13'b111101010110,
13'b111101010111,
13'b111101011010,
13'b111101011011,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101010,
13'b111101101011,
13'b111101101100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111010,
13'b111101111011,
13'b111101111100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001010,
13'b111110001011,
13'b111110001100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011010,
13'b111110011011,
13'b111110011100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101010,
13'b111110101011,
13'b111110101100,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111010,
13'b111110111011,
13'b111111001010,
13'b111111001011,
13'b111111011010,
13'b111111011011,
13'b1000101010110,
13'b1000101010111,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111011,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110001011,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110011011,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110101011,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1001101100101,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110101,
13'b1001110110110,
13'b1010101110101,
13'b1010110000101,
13'b1010110000110,
13'b1010110010101,
13'b1010110010110,
13'b1010110100101,
13'b1010110100110,
13'b1010110110101,
13'b1011110010101,
13'b1011110100101: edge_mask_reg_512p1[77] <= 1'b1;
 		default: edge_mask_reg_512p1[77] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b111000111001,
13'b111000111010,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001001001,
13'b111001001010,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010010100,
13'b1001010010101,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010101,
13'b1100001110101,
13'b1100010000101: edge_mask_reg_512p1[78] <= 1'b1;
 		default: edge_mask_reg_512p1[78] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b1110001010,
13'b10101001100,
13'b10101011011,
13'b10101011100,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11101011011,
13'b11101011100,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001010,
13'b11110001011,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001010,
13'b100110001011,
13'b100110001100,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110001010,
13'b101110001011,
13'b101110001100,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101111010,
13'b110101111011,
13'b110101111100,
13'b110110001010,
13'b110110001011,
13'b110110001100,
13'b110110010111,
13'b110110011000,
13'b110110011010,
13'b110110011011,
13'b110110011100,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110101100,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110110111100,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b111110010111,
13'b111110011000,
13'b111110011010,
13'b111110011011,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110101100,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111110111011,
13'b111110111100,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111001011,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111011011,
13'b111111100111,
13'b111111101000,
13'b1000110010111,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000110111010,
13'b1000110111011,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111001011,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111011011,
13'b1000111100110,
13'b1000111100111,
13'b1001110010111,
13'b1001110100110,
13'b1001110100111,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111100110,
13'b1001111100111,
13'b1010110100110,
13'b1010110100111,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1011110100110,
13'b1011110110101,
13'b1011110110110,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1100110100110,
13'b1100110110110,
13'b1100111000110: edge_mask_reg_512p1[79] <= 1'b1;
 		default: edge_mask_reg_512p1[79] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b1001111000,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111010,
13'b10011111011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b110000111001,
13'b110000111010,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001001,
13'b110011001010,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001001001,
13'b111001001010,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b1000001010110,
13'b1000001010111,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110111,
13'b1000010111000,
13'b1001001010110,
13'b1001001010111,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1010001010110,
13'b1010001010111,
13'b1010001100110,
13'b1010001100111,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110110,
13'b1010010110111,
13'b1011001010110,
13'b1011001100110,
13'b1011001100111,
13'b1011001110101,
13'b1011001110110,
13'b1011001110111,
13'b1011010000101,
13'b1011010000110,
13'b1011010000111,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1100001100110,
13'b1100001100111,
13'b1100001110101,
13'b1100001110110,
13'b1100001110111,
13'b1100010000101,
13'b1100010000110,
13'b1100010000111,
13'b1100010010101,
13'b1100010010110,
13'b1100010010111,
13'b1100010100101,
13'b1100010100110,
13'b1100010100111,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100011000101,
13'b1100011000110,
13'b1101001110101,
13'b1101001110110,
13'b1101001110111,
13'b1101010000101,
13'b1101010000110,
13'b1101010000111,
13'b1101010010101,
13'b1101010010110,
13'b1101010010111,
13'b1101010100101,
13'b1101010100110,
13'b1101010110101,
13'b1101010110110,
13'b1101011000101,
13'b1110001110101,
13'b1110001110110,
13'b1110010000101,
13'b1110010000110,
13'b1110010010101,
13'b1110010010110,
13'b1110010100101,
13'b1110010100110,
13'b1110010110101,
13'b1110010110110,
13'b1111010000110: edge_mask_reg_512p1[80] <= 1'b1;
 		default: edge_mask_reg_512p1[80] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b10001101000,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101001,
13'b100011101010,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b110000111001,
13'b110000111010,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011001,
13'b110011011010,
13'b111001001001,
13'b111001001010,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011001001,
13'b111011001010,
13'b1000001010110,
13'b1000001010111,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100111,
13'b1000010101000,
13'b1000010110111,
13'b1000010111000,
13'b1001001010110,
13'b1001001010111,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010100110,
13'b1001010100111,
13'b1001010110111,
13'b1010001010110,
13'b1010001010111,
13'b1010001100110,
13'b1010001100111,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100110,
13'b1010010100111,
13'b1011001010110,
13'b1011001100110,
13'b1011001100111,
13'b1011001110101,
13'b1011001110110,
13'b1011001110111,
13'b1011010000101,
13'b1011010000110,
13'b1011010000111,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1100001100110,
13'b1100001100111,
13'b1100001110101,
13'b1100001110110,
13'b1100001110111,
13'b1100010000101,
13'b1100010000110,
13'b1100010000111,
13'b1100010010101,
13'b1100010010110,
13'b1100010010111,
13'b1100010100101,
13'b1100010100110,
13'b1100010100111,
13'b1100010110110,
13'b1101001110101,
13'b1101001110110,
13'b1101001110111,
13'b1101010000101,
13'b1101010000110,
13'b1101010000111,
13'b1101010010101,
13'b1101010010110,
13'b1101010010111,
13'b1101010100101,
13'b1101010100110,
13'b1101010100111,
13'b1101010110101,
13'b1101010110110,
13'b1110001110101,
13'b1110001110110,
13'b1110010000101,
13'b1110010000110,
13'b1110010010101,
13'b1110010010110,
13'b1110010100101,
13'b1110010100110,
13'b1110010110110,
13'b1111010000110,
13'b1111010010110,
13'b1111010100110: edge_mask_reg_512p1[81] <= 1'b1;
 		default: edge_mask_reg_512p1[81] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101011001,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101111000,
13'b111101111001,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111101000,
13'b111111101001,
13'b1000110000110,
13'b1000110000111,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010110,
13'b1000111010111,
13'b1001110000110,
13'b1001110000111,
13'b1001110010110,
13'b1001110010111,
13'b1001110100110,
13'b1001110100111,
13'b1001110110110,
13'b1001110110111,
13'b1001111000110,
13'b1001111000111,
13'b1001111010110,
13'b1001111010111,
13'b1010110000110,
13'b1010110000111,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000110,
13'b1010111000111,
13'b1010111010110,
13'b1010111010111,
13'b1010111100110,
13'b1011110000110,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1011110100101,
13'b1011110100110,
13'b1011110100111,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010110,
13'b1011111010111,
13'b1011111100110,
13'b1100110000110,
13'b1100110010101,
13'b1100110010110,
13'b1100110100101,
13'b1100110100110,
13'b1100110110101,
13'b1100110110110,
13'b1100111000101,
13'b1100111000110,
13'b1100111010101,
13'b1100111010110,
13'b1101110010101,
13'b1101110010110,
13'b1101110100101,
13'b1101110100110,
13'b1101110110101,
13'b1101110110110,
13'b1101111000101,
13'b1101111000110,
13'b1101111010101,
13'b1101111010110,
13'b1110110010101,
13'b1110110100101,
13'b1110110100110,
13'b1110110110101,
13'b1110110110110,
13'b1110111000101,
13'b1110111000110,
13'b1110111010101,
13'b1111110010101,
13'b1111110100101,
13'b1111110110101,
13'b1111111000101: edge_mask_reg_512p1[82] <= 1'b1;
 		default: edge_mask_reg_512p1[82] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011001,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000101,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000101,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010100,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b110011111001,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010100,
13'b110110010101,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101000,
13'b110110101001,
13'b111100000100,
13'b111100001001,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001000,
13'b111101001001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011000,
13'b111101011001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101101000,
13'b111101101001,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101111000,
13'b111101111001,
13'b111110000100,
13'b111110000101,
13'b111110001000,
13'b111110001001,
13'b111110010100,
13'b111110010101,
13'b111110011001,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110011,
13'b1000101110100,
13'b1000110000011,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1001101110011,
13'b1001110000011,
13'b1010100100011,
13'b1010100110011,
13'b1010101000011,
13'b1010101010011,
13'b1010101100011: edge_mask_reg_512p1[83] <= 1'b1;
 		default: edge_mask_reg_512p1[83] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001010,
13'b10100001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b110001011001,
13'b110001011010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b1000001110101,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010101,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000100,
13'b1011011000101,
13'b1011011010101,
13'b1100010010100,
13'b1100010010101,
13'b1100010100100,
13'b1100010100101,
13'b1100010110100,
13'b1100010110101,
13'b1100011000100,
13'b1100011000101,
13'b1101010100101,
13'b1101010110101: edge_mask_reg_512p1[84] <= 1'b1;
 		default: edge_mask_reg_512p1[84] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101011,
13'b11010101100,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010011010,
13'b101010011011,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001011100,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001101100,
13'b110001111010,
13'b110001111011,
13'b110010001010,
13'b110010001011,
13'b110010011010,
13'b110010011011,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111000111011,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001001011,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001011011,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001101011,
13'b111001111010,
13'b111001111011,
13'b111010001011,
13'b1000000100111,
13'b1000000101000,
13'b1000000101001,
13'b1000000110111,
13'b1000000111000,
13'b1000000111001,
13'b1000000111010,
13'b1000000111011,
13'b1000001000111,
13'b1000001001000,
13'b1000001001001,
13'b1000001001010,
13'b1000001001011,
13'b1000001010111,
13'b1000001011000,
13'b1000001011001,
13'b1000001011010,
13'b1000001011011,
13'b1000001100111,
13'b1000001101000,
13'b1000001101001,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110110,
13'b1001000110111,
13'b1001000111000,
13'b1001001000110,
13'b1001001000111,
13'b1001001001000,
13'b1001001010111,
13'b1001001011000,
13'b1001001100111,
13'b1001001101000,
13'b1010000010111,
13'b1010000011000,
13'b1010000100110,
13'b1010000100111,
13'b1010000101000,
13'b1010000110110,
13'b1010000110111,
13'b1010000111000,
13'b1010001000110,
13'b1010001000111,
13'b1010001001000,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1010001100111,
13'b1010001101000,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1011000111000,
13'b1011001000110,
13'b1011001000111,
13'b1011001001000,
13'b1011001010110,
13'b1011001010111,
13'b1011001011000,
13'b1011001100111,
13'b1100000010101,
13'b1100000010110,
13'b1100000100101,
13'b1100000100110,
13'b1100000100111,
13'b1100000110101,
13'b1100000110110,
13'b1100000110111,
13'b1100001000110,
13'b1100001000111,
13'b1100001010110,
13'b1100001010111,
13'b1101000010110,
13'b1101000100110,
13'b1101000110110,
13'b1101001000110,
13'b1101001010110: edge_mask_reg_512p1[85] <= 1'b1;
 		default: edge_mask_reg_512p1[85] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100101001,
13'b111100111001,
13'b1000011100011,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1000100100011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[86] <= 1'b1;
 		default: edge_mask_reg_512p1[86] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011001,
13'b11101011010,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b1000011100011,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100100011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011,
13'b1001100100011: edge_mask_reg_512p1[87] <= 1'b1;
 		default: edge_mask_reg_512p1[87] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b1000011100011,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011,
13'b1001100100011: edge_mask_reg_512p1[88] <= 1'b1;
 		default: edge_mask_reg_512p1[88] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1100001010,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101010,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101011000100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1001011110011,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100100011,
13'b1001100110011: edge_mask_reg_512p1[89] <= 1'b1;
 		default: edge_mask_reg_512p1[89] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1100001010,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1001011110011,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100110011: edge_mask_reg_512p1[90] <= 1'b1;
 		default: edge_mask_reg_512p1[90] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100001010,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b100101101010,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b111101001010,
13'b1000011110011,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1010100010011: edge_mask_reg_512p1[91] <= 1'b1;
 		default: edge_mask_reg_512p1[91] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101001,
13'b11101101010,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b100101101010,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b111101001010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011: edge_mask_reg_512p1[92] <= 1'b1;
 		default: edge_mask_reg_512p1[92] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b100101101010,
13'b101011001001,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101001001,
13'b111101001010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101000100,
13'b1001100000011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100: edge_mask_reg_512p1[93] <= 1'b1;
 		default: edge_mask_reg_512p1[93] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100011010,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b100101101010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101000100,
13'b1001100000011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100: edge_mask_reg_512p1[94] <= 1'b1;
 		default: edge_mask_reg_512p1[94] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100011010,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111001,
13'b100101111010,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101000100,
13'b1001100000011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1010100010011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100: edge_mask_reg_512p1[95] <= 1'b1;
 		default: edge_mask_reg_512p1[95] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100101010,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111001,
13'b100101111010,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101010011,
13'b1000101010100,
13'b1001100000011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1010100010011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100: edge_mask_reg_512p1[96] <= 1'b1;
 		default: edge_mask_reg_512p1[96] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100101010,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111001,
13'b11101111010,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111001,
13'b100101111010,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101011001,
13'b111101011010,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101010011,
13'b1000101010100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1010100010011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100: edge_mask_reg_512p1[97] <= 1'b1;
 		default: edge_mask_reg_512p1[97] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100101010,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111001,
13'b100101111010,
13'b101011011001,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101011001,
13'b111101011010,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1010100010011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100: edge_mask_reg_512p1[98] <= 1'b1;
 		default: edge_mask_reg_512p1[98] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100101010,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001010,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111001,
13'b100101111010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b1000100000101,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010100: edge_mask_reg_512p1[99] <= 1'b1;
 		default: edge_mask_reg_512p1[99] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100101010,
13'b1100111010,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001001,
13'b100110001010,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100: edge_mask_reg_512p1[100] <= 1'b1;
 		default: edge_mask_reg_512p1[100] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100111010,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001001,
13'b11110001010,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001001,
13'b100110001010,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100: edge_mask_reg_512p1[101] <= 1'b1;
 		default: edge_mask_reg_512p1[101] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100111010,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001001,
13'b11110001010,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001001,
13'b100110001010,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100: edge_mask_reg_512p1[102] <= 1'b1;
 		default: edge_mask_reg_512p1[102] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100111010,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001001,
13'b100110001010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100100,
13'b1011100110100: edge_mask_reg_512p1[103] <= 1'b1;
 		default: edge_mask_reg_512p1[103] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100111010,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100: edge_mask_reg_512p1[104] <= 1'b1;
 		default: edge_mask_reg_512p1[104] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1101001010,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011001,
13'b100110011010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100: edge_mask_reg_512p1[105] <= 1'b1;
 		default: edge_mask_reg_512p1[105] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1101001010,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011001,
13'b11110011010,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011001,
13'b100110011010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b111100001001,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100: edge_mask_reg_512p1[106] <= 1'b1;
 		default: edge_mask_reg_512p1[106] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1101001010,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011001,
13'b100110011010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100: edge_mask_reg_512p1[107] <= 1'b1;
 		default: edge_mask_reg_512p1[107] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1101001010,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011001,
13'b100110011010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110101,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110101,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[108] <= 1'b1;
 		default: edge_mask_reg_512p1[108] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1101001010,
13'b1101011010,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110101,
13'b1000101110110,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110101,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[109] <= 1'b1;
 		default: edge_mask_reg_512p1[109] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101011010,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110101,
13'b1000101110110,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[110] <= 1'b1;
 		default: edge_mask_reg_512p1[110] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101011010,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101001,
13'b11110101010,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[111] <= 1'b1;
 		default: edge_mask_reg_512p1[111] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101011010,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100001001,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000110,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000101,
13'b1000110000110,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1010101000100,
13'b1010101000101,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101110100,
13'b1100101010100,
13'b1100101100100: edge_mask_reg_512p1[112] <= 1'b1;
 		default: edge_mask_reg_512p1[112] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101011010,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b111110011010,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1010101000100,
13'b1010101000101,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1100101010100,
13'b1100101100100: edge_mask_reg_512p1[113] <= 1'b1;
 		default: edge_mask_reg_512p1[113] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101101010,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b111110011010,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1001110000110,
13'b1010101000100,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1100101100100: edge_mask_reg_512p1[114] <= 1'b1;
 		default: edge_mask_reg_512p1[114] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101101010,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b111110011010,
13'b1000100110101,
13'b1000100110110,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1001100110101,
13'b1001100110110,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1001110000110,
13'b1010101000100,
13'b1010101000101,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1100101100100: edge_mask_reg_512p1[115] <= 1'b1;
 		default: edge_mask_reg_512p1[115] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101101010,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b1000100110101,
13'b1000100110110,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1001100110101,
13'b1001100110110,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1100101100100,
13'b1100101110100: edge_mask_reg_512p1[116] <= 1'b1;
 		default: edge_mask_reg_512p1[116] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b1000011100011,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1010100000011,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1100101010100,
13'b1100101100100,
13'b1100101110100: edge_mask_reg_512p1[117] <= 1'b1;
 		default: edge_mask_reg_512p1[117] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101101010,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b101100011001,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010101,
13'b1010101000101,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1100101100100,
13'b1100101110100: edge_mask_reg_512p1[118] <= 1'b1;
 		default: edge_mask_reg_512p1[118] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100111001,
13'b1000011100011,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100010011: edge_mask_reg_512p1[119] <= 1'b1;
 		default: edge_mask_reg_512p1[119] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100111001,
13'b1000011100011,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[120] <= 1'b1;
 		default: edge_mask_reg_512p1[120] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100111001,
13'b1000011100011,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[121] <= 1'b1;
 		default: edge_mask_reg_512p1[121] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100111001,
13'b1000011100011,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[122] <= 1'b1;
 		default: edge_mask_reg_512p1[122] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[123] <= 1'b1;
 		default: edge_mask_reg_512p1[123] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[124] <= 1'b1;
 		default: edge_mask_reg_512p1[124] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[125] <= 1'b1;
 		default: edge_mask_reg_512p1[125] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[126] <= 1'b1;
 		default: edge_mask_reg_512p1[126] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[127] <= 1'b1;
 		default: edge_mask_reg_512p1[127] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[128] <= 1'b1;
 		default: edge_mask_reg_512p1[128] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[129] <= 1'b1;
 		default: edge_mask_reg_512p1[129] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[130] <= 1'b1;
 		default: edge_mask_reg_512p1[130] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[131] <= 1'b1;
 		default: edge_mask_reg_512p1[131] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[132] <= 1'b1;
 		default: edge_mask_reg_512p1[132] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100: edge_mask_reg_512p1[133] <= 1'b1;
 		default: edge_mask_reg_512p1[133] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100: edge_mask_reg_512p1[134] <= 1'b1;
 		default: edge_mask_reg_512p1[134] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011: edge_mask_reg_512p1[135] <= 1'b1;
 		default: edge_mask_reg_512p1[135] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011110011,
13'b1010100000011,
13'b1010100010011: edge_mask_reg_512p1[136] <= 1'b1;
 		default: edge_mask_reg_512p1[136] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011110011,
13'b1010100000011,
13'b1010100010011: edge_mask_reg_512p1[137] <= 1'b1;
 		default: edge_mask_reg_512p1[137] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011110011,
13'b1010100000011,
13'b1010100010011: edge_mask_reg_512p1[138] <= 1'b1;
 		default: edge_mask_reg_512p1[138] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011110011,
13'b1010100000011,
13'b1010100010011: edge_mask_reg_512p1[139] <= 1'b1;
 		default: edge_mask_reg_512p1[139] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011110011,
13'b1010100000011,
13'b1010100010011: edge_mask_reg_512p1[140] <= 1'b1;
 		default: edge_mask_reg_512p1[140] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011110011,
13'b1010100000011,
13'b1010100010011: edge_mask_reg_512p1[141] <= 1'b1;
 		default: edge_mask_reg_512p1[141] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010100000011,
13'b1010100010011: edge_mask_reg_512p1[142] <= 1'b1;
 		default: edge_mask_reg_512p1[142] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[143] <= 1'b1;
 		default: edge_mask_reg_512p1[143] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[144] <= 1'b1;
 		default: edge_mask_reg_512p1[144] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[145] <= 1'b1;
 		default: edge_mask_reg_512p1[145] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[146] <= 1'b1;
 		default: edge_mask_reg_512p1[146] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[147] <= 1'b1;
 		default: edge_mask_reg_512p1[147] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[148] <= 1'b1;
 		default: edge_mask_reg_512p1[148] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[149] <= 1'b1;
 		default: edge_mask_reg_512p1[149] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010110100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011000100,
13'b111011001001,
13'b111011001010,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100110100,
13'b111100111001,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[150] <= 1'b1;
 		default: edge_mask_reg_512p1[150] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010110,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100111001,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[151] <= 1'b1;
 		default: edge_mask_reg_512p1[151] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010110100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010010,
13'b111011010011,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100111001,
13'b1000011010011,
13'b1000011100011,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[152] <= 1'b1;
 		default: edge_mask_reg_512p1[152] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010110100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b1000011010011,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[153] <= 1'b1;
 		default: edge_mask_reg_512p1[153] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011111010,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001001,
13'b11101001010,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100111001,
13'b110100111010,
13'b111011001001,
13'b111011001010,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011011001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b1000011010011,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1001011010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[154] <= 1'b1;
 		default: edge_mask_reg_512p1[154] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011111010,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001001,
13'b11101001010,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010110100,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111010111001,
13'b111011001001,
13'b111011001010,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1001011010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011: edge_mask_reg_512p1[155] <= 1'b1;
 		default: edge_mask_reg_512p1[155] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011101010,
13'b1011111010,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b110010101001,
13'b110010110100,
13'b110010110101,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1001011010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011: edge_mask_reg_512p1[156] <= 1'b1;
 		default: edge_mask_reg_512p1[156] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011101010,
13'b1011111010,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001010,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111001,
13'b100100111010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111010110100,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b1000011000011,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1001011010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011: edge_mask_reg_512p1[157] <= 1'b1;
 		default: edge_mask_reg_512p1[157] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011101010,
13'b1011111001,
13'b1011111010,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b1000011000011,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001100000011: edge_mask_reg_512p1[158] <= 1'b1;
 		default: edge_mask_reg_512p1[158] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011101010,
13'b1011111001,
13'b1011111010,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111001,
13'b11100111010,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b1000011000011,
13'b1000011000100,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1001011000011,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1010011010011: edge_mask_reg_512p1[159] <= 1'b1;
 		default: edge_mask_reg_512p1[159] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011101010,
13'b1011111001,
13'b1011111010,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010100100,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b1000011000011,
13'b1000011000100,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1010011010011: edge_mask_reg_512p1[160] <= 1'b1;
 		default: edge_mask_reg_512p1[160] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011011010,
13'b1011101010,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010100100,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b1000011000011,
13'b1000011000100,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1010011000011,
13'b1010011010011,
13'b1010011100011,
13'b1010011110011: edge_mask_reg_512p1[161] <= 1'b1;
 		default: edge_mask_reg_512p1[161] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011011010,
13'b1011101010,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100101,
13'b11010100110,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101001,
13'b100100101010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010100100,
13'b111010100101,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b1000010110011,
13'b1000011000011,
13'b1000011000100,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011110011: edge_mask_reg_512p1[162] <= 1'b1;
 		default: edge_mask_reg_512p1[162] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011011010,
13'b1011101001,
13'b1011101010,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101001,
13'b100100101010,
13'b101010001001,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010100100,
13'b111010100101,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b1000010110011,
13'b1000010110100,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1001010110011,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011: edge_mask_reg_512p1[163] <= 1'b1;
 		default: edge_mask_reg_512p1[163] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011011010,
13'b1011101001,
13'b1011101010,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101001,
13'b11100101010,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101001,
13'b100100101010,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b111010011001,
13'b111010100100,
13'b111010100101,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1001010110011,
13'b1001010110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100: edge_mask_reg_512p1[164] <= 1'b1;
 		default: edge_mask_reg_512p1[164] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011011010,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101001,
13'b100100101010,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100001001,
13'b111100001010,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1001010110011,
13'b1001010110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100: edge_mask_reg_512p1[165] <= 1'b1;
 		default: edge_mask_reg_512p1[165] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1011001010,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101001,
13'b101010001001,
13'b101010001010,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b111010010100,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100001001,
13'b111100001010,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1001010110011,
13'b1001010110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100: edge_mask_reg_512p1[166] <= 1'b1;
 		default: edge_mask_reg_512p1[166] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1011001010,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011001,
13'b100100011010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b111010010100,
13'b111010010101,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1001010100011,
13'b1001010110011,
13'b1001010110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100: edge_mask_reg_512p1[167] <= 1'b1;
 		default: edge_mask_reg_512p1[167] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1011001010,
13'b1011011001,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011001,
13'b11100011010,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011001,
13'b100100011010,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b111010010100,
13'b111010010101,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1001010100011,
13'b1001010100100,
13'b1001010110011,
13'b1001010110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1011010110100: edge_mask_reg_512p1[168] <= 1'b1;
 		default: edge_mask_reg_512p1[168] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1011001010,
13'b1011011001,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011001,
13'b11100011010,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011001,
13'b100100011010,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1001010100011,
13'b1001010100100,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1011010110100: edge_mask_reg_512p1[169] <= 1'b1;
 		default: edge_mask_reg_512p1[169] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1011001010,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011001,
13'b100100011010,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b110001111001,
13'b110001111010,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011111001,
13'b111011111010,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1001010100011,
13'b1001010100100,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[170] <= 1'b1;
 		default: edge_mask_reg_512p1[170] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010111010,
13'b1011001010,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001001,
13'b100100001010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b110001111001,
13'b110001111010,
13'b110010000110,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[171] <= 1'b1;
 		default: edge_mask_reg_512p1[171] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010111010,
13'b1011001001,
13'b1011001010,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001001,
13'b100100001010,
13'b101001101001,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b111010000100,
13'b111010000101,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010100,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1001010010011,
13'b1001010010100,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010100,
13'b1010010010011,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[172] <= 1'b1;
 		default: edge_mask_reg_512p1[172] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010111010,
13'b1011001001,
13'b1011001010,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001001,
13'b11100001010,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001001,
13'b100100001010,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111010000100,
13'b111010000101,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b1000010000101,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010100,
13'b1001011010101,
13'b1010010010011,
13'b1010010010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[173] <= 1'b1;
 		default: edge_mask_reg_512p1[173] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010111010,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001001,
13'b100100001010,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b1000010000100,
13'b1000010000101,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1001010000101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010101,
13'b1010010010011,
13'b1010010010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[174] <= 1'b1;
 		default: edge_mask_reg_512p1[174] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010111010,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001001,
13'b100100001010,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001101001,
13'b110001101010,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011101001,
13'b111011101010,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1001010000101,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010101,
13'b1010010010011,
13'b1010010010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000011,
13'b1010011000100,
13'b1011010010100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[175] <= 1'b1;
 		default: edge_mask_reg_512p1[175] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001010,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001101001,
13'b110001101010,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011101001,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1001010000101,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011010101,
13'b1010010010100,
13'b1010010010101,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000100,
13'b1011010010100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[176] <= 1'b1;
 		default: edge_mask_reg_512p1[176] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010111001,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001011001,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001101001,
13'b110001101010,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1001010000100,
13'b1001010000101,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011010101,
13'b1010010000100,
13'b1010010010100,
13'b1010010010101,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000100,
13'b1011010010100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[177] <= 1'b1;
 		default: edge_mask_reg_512p1[177] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011010,
13'b1010101010,
13'b1010111001,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111001,
13'b11011111010,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001101001,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b1000001110101,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000101,
13'b1001011000110,
13'b1010010000100,
13'b1010010010100,
13'b1010010010101,
13'b1010010100100,
13'b1010010100101,
13'b1010010110100,
13'b1010010110101,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010110100,
13'b1100010010100: edge_mask_reg_512p1[178] <= 1'b1;
 		default: edge_mask_reg_512p1[178] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011010,
13'b1010101010,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111010,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000101,
13'b1001011000110,
13'b1010010000100,
13'b1010010010100,
13'b1010010010101,
13'b1010010100100,
13'b1010010100101,
13'b1010010110100,
13'b1010010110101,
13'b1011010000100,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1100010010100: edge_mask_reg_512p1[179] <= 1'b1;
 		default: edge_mask_reg_512p1[179] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b1001111000,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011010,
13'b1010101010,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b110001011001,
13'b110001011010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000101,
13'b1001011000110,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1010010100100,
13'b1010010100101,
13'b1010010110100,
13'b1010010110101,
13'b1011010000100,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1100010010100: edge_mask_reg_512p1[180] <= 1'b1;
 		default: edge_mask_reg_512p1[180] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b1001111000,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011010,
13'b1010101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101001,
13'b100011101010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b110001011001,
13'b110001011010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000101,
13'b1001011000110,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1010010100100,
13'b1010010100101,
13'b1010010110100,
13'b1010010110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1100010010100: edge_mask_reg_512p1[181] <= 1'b1;
 		default: edge_mask_reg_512p1[181] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001010,
13'b1001111000,
13'b1001111001,
13'b1010001010,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b10001101000,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101001,
13'b11011101010,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101001,
13'b100011101010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b110001011001,
13'b110001011010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001100110,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110101,
13'b1001010110110,
13'b1001011000101,
13'b1010001110100,
13'b1010001110101,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1011001110100,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1100010000100,
13'b1100010010100: edge_mask_reg_512p1[182] <= 1'b1;
 		default: edge_mask_reg_512p1[182] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011010,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110001011001,
13'b110001011010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111001100110,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1010001110100,
13'b1010001110101,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1011001110100,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1011011000100,
13'b1011011010100,
13'b1100010000100,
13'b1100010010100,
13'b1100010100100: edge_mask_reg_512p1[183] <= 1'b1;
 		default: edge_mask_reg_512p1[183] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001010,
13'b1001111000,
13'b1001111001,
13'b1010001010,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b11001011000,
13'b11001011001,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101001,
13'b11011101010,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101001,
13'b100011101010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100110,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100110,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011001,
13'b110011011010,
13'b111001100101,
13'b111001100110,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011001001,
13'b111011001010,
13'b1000001100101,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110101,
13'b1000010110110,
13'b1001001100101,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110101,
13'b1001010110110,
13'b1010001110100,
13'b1010001110101,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110101,
13'b1011001110100,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1100010000100,
13'b1100010010100: edge_mask_reg_512p1[184] <= 1'b1;
 		default: edge_mask_reg_512p1[184] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[185] <= 1'b1;
 		default: edge_mask_reg_512p1[185] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011010,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1001011100011,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011: edge_mask_reg_512p1[186] <= 1'b1;
 		default: edge_mask_reg_512p1[186] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011001,
13'b11101011010,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010100: edge_mask_reg_512p1[187] <= 1'b1;
 		default: edge_mask_reg_512p1[187] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010100,
13'b1010100100100: edge_mask_reg_512p1[188] <= 1'b1;
 		default: edge_mask_reg_512p1[188] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1100001010,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101010,
13'b10101101011,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010100,
13'b1010100100100: edge_mask_reg_512p1[189] <= 1'b1;
 		default: edge_mask_reg_512p1[189] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101010,
13'b10101101011,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101011001001,
13'b101011001010,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b111101001010,
13'b1000011100100,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1001100100100,
13'b1001100110100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100100,
13'b1010100110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[190] <= 1'b1;
 		default: edge_mask_reg_512p1[190] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b100101101010,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b101101101010,
13'b110011001001,
13'b110011001010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100011,
13'b1010100100100,
13'b1010100110100,
13'b1011100000100,
13'b1011100010100,
13'b1011100100100: edge_mask_reg_512p1[191] <= 1'b1;
 		default: edge_mask_reg_512p1[191] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101010,
13'b11101101011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1001011110100,
13'b1001011110101,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1001100110101,
13'b1010100000100,
13'b1010100010100,
13'b1010100010101,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1011100000100,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100: edge_mask_reg_512p1[192] <= 1'b1;
 		default: edge_mask_reg_512p1[192] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011100110,
13'b110011100111,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b1000011100101,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1001011110101,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1001100110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1010100110101,
13'b1011100000100,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1100100100101: edge_mask_reg_512p1[193] <= 1'b1;
 		default: edge_mask_reg_512p1[193] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1010100110101,
13'b1010101000100,
13'b1011100000100,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1100100100101: edge_mask_reg_512p1[194] <= 1'b1;
 		default: edge_mask_reg_512p1[194] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b110011110110,
13'b110011110111,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b1000011110101,
13'b1000011110110,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110101,
13'b1000100110110,
13'b1001011110101,
13'b1001011110110,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1010100110101,
13'b1010101000100,
13'b1010101000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1011101000101,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100110101: edge_mask_reg_512p1[195] <= 1'b1;
 		default: edge_mask_reg_512p1[195] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100011001010,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b110011110110,
13'b110011110111,
13'b110011111001,
13'b110011111010,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000011110101,
13'b1000011110110,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110101,
13'b1000100110110,
13'b1001011110110,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000101,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010101000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1011101000101,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100110101: edge_mask_reg_512p1[196] <= 1'b1;
 		default: edge_mask_reg_512p1[196] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111010,
13'b11101111011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111010,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110101,
13'b1000100110110,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110101,
13'b1001100110110,
13'b1001101000101,
13'b1010100000101,
13'b1010100000110,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010101000101,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011101000101,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100110101,
13'b1100101000101: edge_mask_reg_512p1[197] <= 1'b1;
 		default: edge_mask_reg_512p1[197] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111010,
13'b11101111011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000101,
13'b1010100000101,
13'b1010100000110,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010101000101,
13'b1011100010101,
13'b1011100010110,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011101000101,
13'b1100100100101,
13'b1100100110101,
13'b1100101000101: edge_mask_reg_512p1[198] <= 1'b1;
 		default: edge_mask_reg_512p1[198] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111010,
13'b11101111011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000101,
13'b1001101000110,
13'b1010100000110,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000101,
13'b1010101000110,
13'b1011100010101,
13'b1011100010110,
13'b1011100100101,
13'b1011100100110,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011101000101,
13'b1011101000110,
13'b1100100100101,
13'b1100100110101,
13'b1100100110110,
13'b1100101000101,
13'b1100101000110,
13'b1101100100101,
13'b1101100110101,
13'b1101101000101: edge_mask_reg_512p1[199] <= 1'b1;
 		default: edge_mask_reg_512p1[199] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001010,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111010,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000100000101,
13'b1000100000110,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1001100000110,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000101,
13'b1001101000110,
13'b1010100000110,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000101,
13'b1010101000110,
13'b1011100010110,
13'b1011100100101,
13'b1011100100110,
13'b1011100110101,
13'b1011100110110,
13'b1011101000101,
13'b1011101000110,
13'b1011101010101,
13'b1100100100101,
13'b1100100100110,
13'b1100100110101,
13'b1100100110110,
13'b1100101000101,
13'b1100101000110,
13'b1101100100101,
13'b1101100110101,
13'b1101101000101,
13'b1101101000110: edge_mask_reg_512p1[200] <= 1'b1;
 		default: edge_mask_reg_512p1[200] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001010,
13'b10110001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b111101101010,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000101,
13'b1001101000110,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000101,
13'b1010101000110,
13'b1011100010110,
13'b1011100010111,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101010101,
13'b1100100100101,
13'b1100100100110,
13'b1100100110101,
13'b1100100110110,
13'b1100101000101,
13'b1100101000110,
13'b1100101010101,
13'b1101100100101,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110: edge_mask_reg_512p1[201] <= 1'b1;
 		default: edge_mask_reg_512p1[201] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001010,
13'b10110001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1011100010110,
13'b1011100010111,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1100100100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101010101,
13'b1100101010110,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010110: edge_mask_reg_512p1[202] <= 1'b1;
 		default: edge_mask_reg_512p1[202] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001010,
13'b10110001011,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001010,
13'b11110001011,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001010,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1011100010110,
13'b1011100010111,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101010101,
13'b1100101010110,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010110,
13'b1110100110110: edge_mask_reg_512p1[203] <= 1'b1;
 		default: edge_mask_reg_512p1[203] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111010,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1011100010110,
13'b1011100010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010110,
13'b1110100110110,
13'b1110101000110: edge_mask_reg_512p1[204] <= 1'b1;
 		default: edge_mask_reg_512p1[204] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010110,
13'b1000100010111,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111010,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101011000,
13'b1001100010110,
13'b1001100010111,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010111,
13'b1001101011000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1011100010110,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010110,
13'b1110100110110,
13'b1110101000110: edge_mask_reg_512p1[205] <= 1'b1;
 		default: edge_mask_reg_512p1[205] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001010,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101001010,
13'b1000101010111,
13'b1000101011000,
13'b1001100010110,
13'b1001100010111,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010111,
13'b1001101011000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010111,
13'b1011100010110,
13'b1011100010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010110,
13'b1110101000110,
13'b1110101010110: edge_mask_reg_512p1[206] <= 1'b1;
 		default: edge_mask_reg_512p1[206] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001010,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b111101111010,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101010111,
13'b1000101011000,
13'b1001100010110,
13'b1001100010111,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010111,
13'b1001101011000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1010100100111,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010111,
13'b1010101011000,
13'b1011100010110,
13'b1011100010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1100100100110,
13'b1100100100111,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101010110,
13'b1110101000110,
13'b1110101010110: edge_mask_reg_512p1[207] <= 1'b1;
 		default: edge_mask_reg_512p1[207] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011011,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b111100001001,
13'b111100001010,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101001,
13'b111101101010,
13'b111101111010,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101010111,
13'b1000101011000,
13'b1001100010111,
13'b1001100011000,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1010100100111,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010111,
13'b1010101011000,
13'b1011100010110,
13'b1011100010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1100100100110,
13'b1100100100111,
13'b1100100110110,
13'b1100100110111,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1101100110110,
13'b1101100110111,
13'b1101101000110,
13'b1101101000111,
13'b1101101010110,
13'b1110101000110,
13'b1110101010110: edge_mask_reg_512p1[208] <= 1'b1;
 		default: edge_mask_reg_512p1[208] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011010,
13'b11110011011,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b111100001001,
13'b111100001010,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101010,
13'b111101111010,
13'b1000100010111,
13'b1000100011000,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101010111,
13'b1000101011000,
13'b1001100010111,
13'b1001100011000,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1010100010111,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010111,
13'b1010101011000,
13'b1011100010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1100100100111,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1101100110110,
13'b1101100110111,
13'b1101101000110,
13'b1101101000111,
13'b1101101010110,
13'b1101101010111,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110: edge_mask_reg_512p1[209] <= 1'b1;
 		default: edge_mask_reg_512p1[209] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011010,
13'b11110011011,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101010,
13'b111101111010,
13'b1000100011000,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1001100011000,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101101000,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010111,
13'b1010101011000,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1100100100111,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1101100110110,
13'b1101100110111,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1111101000110,
13'b1111101010110: edge_mask_reg_512p1[210] <= 1'b1;
 		default: edge_mask_reg_512p1[210] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011010,
13'b11110011011,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b100110011011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110011011,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b111100001010,
13'b111100001011,
13'b111100011010,
13'b111100011011,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101010,
13'b111101101011,
13'b111101111010,
13'b111101111011,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1001100100111,
13'b1001100101000,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1010100100111,
13'b1010100101000,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101101000,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1100100100111,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111: edge_mask_reg_512p1[211] <= 1'b1;
 		default: edge_mask_reg_512p1[211] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011010,
13'b11110011011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b100110011011,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110011011,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011010,
13'b111100001010,
13'b111100001011,
13'b111100011010,
13'b111100011011,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111010,
13'b111101111011,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1001100100111,
13'b1001100101000,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1010100100111,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1011100100111,
13'b1011100101000,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1011101101000,
13'b1100100100111,
13'b1100100101000,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1100101101000,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1110101100110,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111: edge_mask_reg_512p1[212] <= 1'b1;
 		default: edge_mask_reg_512p1[212] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b100110011011,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110011011,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011010,
13'b110110011011,
13'b111100001010,
13'b111100001011,
13'b111100011010,
13'b111100011011,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1010100100111,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1011100100111,
13'b1011100101000,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1011101101000,
13'b1100100100111,
13'b1100100101000,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1100101101000,
13'b1101100100111,
13'b1101100101000,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1110101100110,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111: edge_mask_reg_512p1[213] <= 1'b1;
 		default: edge_mask_reg_512p1[213] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b100110011011,
13'b100110101010,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110011011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011010,
13'b110110011011,
13'b111100001010,
13'b111100001011,
13'b111100011010,
13'b111100011011,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b1000100101000,
13'b1000100101001,
13'b1000100111000,
13'b1000100111001,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1000101101001,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101001000,
13'b1001101001001,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1001101101001,
13'b1010100100111,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1011100100111,
13'b1011100101000,
13'b1011100110111,
13'b1011100111000,
13'b1011101000111,
13'b1011101001000,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1011101101000,
13'b1100100100111,
13'b1100100101000,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1100101101000,
13'b1101100100111,
13'b1101100101000,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1110101100110,
13'b1110101100111,
13'b1111101000111,
13'b1111101010111: edge_mask_reg_512p1[214] <= 1'b1;
 		default: edge_mask_reg_512p1[214] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101010,
13'b100110101011,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110011011,
13'b101110101010,
13'b101110101011,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011010,
13'b110110011011,
13'b111100001010,
13'b111100011010,
13'b111100011011,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b1000100111000,
13'b1000100111001,
13'b1000101001000,
13'b1000101001001,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1000101101001,
13'b1001100101000,
13'b1001100101001,
13'b1001100111000,
13'b1001100111001,
13'b1001101001000,
13'b1001101001001,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1001101101001,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101101000,
13'b1010101101001,
13'b1011100101000,
13'b1011100110111,
13'b1011100111000,
13'b1011100111001,
13'b1011101000111,
13'b1011101001000,
13'b1011101010111,
13'b1011101011000,
13'b1011101011001,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1100100101000,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1100101101000,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100111,
13'b1101101101000,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100111,
13'b1111101000111,
13'b1111101010111: edge_mask_reg_512p1[215] <= 1'b1;
 		default: edge_mask_reg_512p1[215] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101010,
13'b100110101011,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110011011,
13'b101110101010,
13'b101110101011,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011010,
13'b110110011011,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000101,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1000101101001,
13'b1001011100011,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1001101101001,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1011100000100,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011100111001,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101011001,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1100101101000,
13'b1101100100101,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1110100110110,
13'b1110100110111,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111: edge_mask_reg_512p1[216] <= 1'b1;
 		default: edge_mask_reg_512p1[216] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101010,
13'b100110101011,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101010,
13'b101110101011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110110,
13'b1010101110111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011100111001,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101011001,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100101,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000100,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010100,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100100,
13'b1101101100101,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1110100110101,
13'b1110101000100,
13'b1110101000101,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101010100,
13'b1110101010101,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100100,
13'b1110101100101,
13'b1110101100110,
13'b1110101100111,
13'b1111101000101,
13'b1111101000110,
13'b1111101000111,
13'b1111101010101,
13'b1111101010110,
13'b1111101010111: edge_mask_reg_512p1[217] <= 1'b1;
 		default: edge_mask_reg_512p1[217] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b1000011100011,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[218] <= 1'b1;
 		default: edge_mask_reg_512p1[218] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[219] <= 1'b1;
 		default: edge_mask_reg_512p1[219] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[220] <= 1'b1;
 		default: edge_mask_reg_512p1[220] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100: edge_mask_reg_512p1[221] <= 1'b1;
 		default: edge_mask_reg_512p1[221] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011110011,
13'b1010100000011,
13'b1010100010011: edge_mask_reg_512p1[222] <= 1'b1;
 		default: edge_mask_reg_512p1[222] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[223] <= 1'b1;
 		default: edge_mask_reg_512p1[223] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[224] <= 1'b1;
 		default: edge_mask_reg_512p1[224] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[225] <= 1'b1;
 		default: edge_mask_reg_512p1[225] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[226] <= 1'b1;
 		default: edge_mask_reg_512p1[226] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100: edge_mask_reg_512p1[227] <= 1'b1;
 		default: edge_mask_reg_512p1[227] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1010011100100,
13'b1010011110100,
13'b1010100000100,
13'b1010100010100,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[228] <= 1'b1;
 		default: edge_mask_reg_512p1[228] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100101,
13'b1000100100110,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100010100,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[229] <= 1'b1;
 		default: edge_mask_reg_512p1[229] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100101,
13'b1000100100110,
13'b1001011010101,
13'b1001011100100,
13'b1001011100101,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100100101,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[230] <= 1'b1;
 		default: edge_mask_reg_512p1[230] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100101,
13'b1000100100110,
13'b1001011010101,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[231] <= 1'b1;
 		default: edge_mask_reg_512p1[231] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011011001,
13'b110011011010,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100101,
13'b1000100100110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011011100100,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101: edge_mask_reg_512p1[232] <= 1'b1;
 		default: edge_mask_reg_512p1[232] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011011001,
13'b110011011010,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100101,
13'b1000100100110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011011100100,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1100011110100,
13'b1100100000100: edge_mask_reg_512p1[233] <= 1'b1;
 		default: edge_mask_reg_512p1[233] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011001,
13'b110011011010,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1011011100100,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000100,
13'b1100100000101: edge_mask_reg_512p1[234] <= 1'b1;
 		default: edge_mask_reg_512p1[234] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011010110,
13'b110011010111,
13'b110011011001,
13'b110011011010,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011010110,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100101,
13'b1010100100110,
13'b1011011100100,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1100011110100,
13'b1100011110101,
13'b1100100000100,
13'b1100100000101: edge_mask_reg_512p1[235] <= 1'b1;
 		default: edge_mask_reg_512p1[235] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011010110,
13'b110011010111,
13'b110011011001,
13'b110011011010,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011010110,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100101,
13'b1010100100110,
13'b1011011100100,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1100011110100,
13'b1100011110101,
13'b1100100000100,
13'b1100100000101: edge_mask_reg_512p1[236] <= 1'b1;
 		default: edge_mask_reg_512p1[236] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011010110,
13'b110011010111,
13'b110011011001,
13'b110011011010,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011010110,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100101,
13'b1010100100110,
13'b1011011100100,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1100011110101,
13'b1100100000101: edge_mask_reg_512p1[237] <= 1'b1;
 		default: edge_mask_reg_512p1[237] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100111,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011010110,
13'b110011010111,
13'b110011011001,
13'b110011011010,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1001011010101,
13'b1001011010110,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001100000101,
13'b1001100000110,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100101,
13'b1010100100110,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100010100,
13'b1100011110101,
13'b1100100000101: edge_mask_reg_512p1[238] <= 1'b1;
 		default: edge_mask_reg_512p1[238] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011010110,
13'b110011010111,
13'b110011011001,
13'b110011011010,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1001011010101,
13'b1001011010110,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001100000101,
13'b1001100000110,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010101,
13'b1010100010110,
13'b1010100100101,
13'b1010100100110,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1100011110101,
13'b1100100000101: edge_mask_reg_512p1[239] <= 1'b1;
 		default: edge_mask_reg_512p1[239] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011010110,
13'b110011010111,
13'b110011011001,
13'b110011011010,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100110,
13'b1000100100111,
13'b1001011010110,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100100110,
13'b1011011100101,
13'b1011011100110,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100010101,
13'b1011100010110,
13'b1100011110101,
13'b1100100000101,
13'b1101011110101,
13'b1101100000101: edge_mask_reg_512p1[240] <= 1'b1;
 		default: edge_mask_reg_512p1[240] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1001011010110,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100110,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1011011100101,
13'b1011011100110,
13'b1011011110101,
13'b1011011110110,
13'b1011100000101,
13'b1011100000110,
13'b1011100010101,
13'b1011100010110,
13'b1100011110101,
13'b1100011110110,
13'b1100100000101,
13'b1100100000110,
13'b1101011110101,
13'b1101100000101: edge_mask_reg_512p1[241] <= 1'b1;
 		default: edge_mask_reg_512p1[241] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010110,
13'b1000011010111,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1001011010110,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010110,
13'b1001100010111,
13'b1001100100110,
13'b1001100100111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1011011100101,
13'b1011011100110,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010101,
13'b1011100010110,
13'b1100011110101,
13'b1100011110110,
13'b1100100000101,
13'b1100100000110,
13'b1101011110101,
13'b1101100000101: edge_mask_reg_512p1[242] <= 1'b1;
 		default: edge_mask_reg_512p1[242] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010111,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010110,
13'b1001100010111,
13'b1001100100110,
13'b1001100100111,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010110,
13'b1011100010111,
13'b1100011110101,
13'b1100011110110,
13'b1100100000101,
13'b1100100000110,
13'b1101011110101,
13'b1101100000101: edge_mask_reg_512p1[243] <= 1'b1;
 		default: edge_mask_reg_512p1[243] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010111,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1001011010111,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010110,
13'b1001100010111,
13'b1001100100110,
13'b1001100100111,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010110,
13'b1011100010111,
13'b1100011110101,
13'b1100011110110,
13'b1100100000101,
13'b1100100000110,
13'b1101011110101,
13'b1101011110110,
13'b1101100000101,
13'b1101100000110: edge_mask_reg_512p1[244] <= 1'b1;
 		default: edge_mask_reg_512p1[244] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011010,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010111,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1001011010111,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100110,
13'b1001100100111,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010110,
13'b1011100010111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1101011110101,
13'b1101011110110,
13'b1101100000101,
13'b1101100000110: edge_mask_reg_512p1[245] <= 1'b1;
 		default: edge_mask_reg_512p1[245] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011010,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1001011010111,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100110,
13'b1001100100111,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010110,
13'b1010100010111,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010110,
13'b1011100010111,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1101011110101,
13'b1101011110110,
13'b1101100000101,
13'b1101100000110: edge_mask_reg_512p1[246] <= 1'b1;
 		default: edge_mask_reg_512p1[246] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011010,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110111,
13'b1000011111000,
13'b1000100000111,
13'b1000100001000,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1001011010111,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1010011100110,
13'b1010011100111,
13'b1010011110110,
13'b1010011110111,
13'b1010100000110,
13'b1010100000111,
13'b1010100010110,
13'b1010100010111,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010110,
13'b1011100010111,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1101011110101,
13'b1101011110110,
13'b1101100000101,
13'b1101100000110,
13'b1110011110110,
13'b1110100000110: edge_mask_reg_512p1[247] <= 1'b1;
 		default: edge_mask_reg_512p1[247] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011010,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100111,
13'b1000011101000,
13'b1000011110111,
13'b1000011111000,
13'b1000100000111,
13'b1000100001000,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1001011010111,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110110,
13'b1010011110111,
13'b1010100000110,
13'b1010100000111,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010110,
13'b1011100010111,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1101011110101,
13'b1101011110110,
13'b1101100000101,
13'b1101100000110,
13'b1110011110110,
13'b1110100000110: edge_mask_reg_512p1[248] <= 1'b1;
 		default: edge_mask_reg_512p1[248] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110100,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011010,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100101,
13'b1001100100110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1010100100101,
13'b1010100100110,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010100,
13'b1011100010110,
13'b1011100010111,
13'b1100011100110,
13'b1100011100111,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1101011110101,
13'b1101011110110,
13'b1101100000101,
13'b1101100000110,
13'b1110011110110,
13'b1110100000110: edge_mask_reg_512p1[249] <= 1'b1;
 		default: edge_mask_reg_512p1[249] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011010,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100101,
13'b1001100100110,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1010100100101,
13'b1010100100110,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100100101,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010101,
13'b1100100010110,
13'b1100100010111,
13'b1101011110100,
13'b1101011110101,
13'b1101011110110,
13'b1101100000100,
13'b1101100000101,
13'b1101100000110,
13'b1110011110100,
13'b1110011110101,
13'b1110011110110,
13'b1110100000100,
13'b1110100000101,
13'b1110100000110: edge_mask_reg_512p1[250] <= 1'b1;
 		default: edge_mask_reg_512p1[250] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[251] <= 1'b1;
 		default: edge_mask_reg_512p1[251] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011000100,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011: edge_mask_reg_512p1[252] <= 1'b1;
 		default: edge_mask_reg_512p1[252] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011000100,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b1000011010011,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000100: edge_mask_reg_512p1[253] <= 1'b1;
 		default: edge_mask_reg_512p1[253] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011111010,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001001,
13'b11101001010,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000100,
13'b1010100010100: edge_mask_reg_512p1[254] <= 1'b1;
 		default: edge_mask_reg_512p1[254] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011111010,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100101001,
13'b111100101010,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000100,
13'b1010100010100: edge_mask_reg_512p1[255] <= 1'b1;
 		default: edge_mask_reg_512p1[255] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b1000011000101,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010100,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000100,
13'b1010100010100,
13'b1011011110100: edge_mask_reg_512p1[256] <= 1'b1;
 		default: edge_mask_reg_512p1[256] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010101001,
13'b110010101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b1000011000101,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010100,
13'b1001011010100,
13'b1001011010101,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100010100,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100: edge_mask_reg_512p1[257] <= 1'b1;
 		default: edge_mask_reg_512p1[257] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001010,
13'b10101001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010101001,
13'b110010101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100010100,
13'b1001011000101,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010100,
13'b1010011010100,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1011011100100,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100: edge_mask_reg_512p1[258] <= 1'b1;
 		default: edge_mask_reg_512p1[258] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001010,
13'b10101001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1001011000101,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100010100,
13'b1010011010100,
13'b1010011010101,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101: edge_mask_reg_512p1[259] <= 1'b1;
 		default: edge_mask_reg_512p1[259] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001010,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b110100111010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1001011000101,
13'b1001011000110,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110101: edge_mask_reg_512p1[260] <= 1'b1;
 		default: edge_mask_reg_512p1[260] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000101,
13'b1000100000110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1010011000101,
13'b1010011000110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110101,
13'b1100100000101: edge_mask_reg_512p1[261] <= 1'b1;
 		default: edge_mask_reg_512p1[261] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111010,
13'b11100111011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000100000101,
13'b1000100000110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000101,
13'b1010011000101,
13'b1010011000110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110101,
13'b1100100000101: edge_mask_reg_512p1[262] <= 1'b1;
 		default: edge_mask_reg_512p1[262] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111010,
13'b11100111011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111010,
13'b110010011001,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000100000101,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001100000101,
13'b1010011000101,
13'b1010011000110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1100011100101,
13'b1100011110101,
13'b1100100000101: edge_mask_reg_512p1[263] <= 1'b1;
 		default: edge_mask_reg_512p1[263] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001011,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b110010011001,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001100000101,
13'b1010011000101,
13'b1010011000110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100101,
13'b1010011100110,
13'b1010011110101,
13'b1010011110110,
13'b1010100000101,
13'b1011011010101,
13'b1011011010110,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000101,
13'b1100011010101,
13'b1100011100101,
13'b1100011110101,
13'b1100100000101,
13'b1101011100101: edge_mask_reg_512p1[264] <= 1'b1;
 		default: edge_mask_reg_512p1[264] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001011,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b101010001010,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110101,
13'b1000011110110,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010100000101,
13'b1011011000110,
13'b1011011010101,
13'b1011011010110,
13'b1011011100101,
13'b1011011100110,
13'b1011011110101,
13'b1011011110110,
13'b1011100000101,
13'b1100011010101,
13'b1100011010110,
13'b1100011100101,
13'b1100011110101,
13'b1100100000101,
13'b1101011100101,
13'b1101011110101: edge_mask_reg_512p1[265] <= 1'b1;
 		default: edge_mask_reg_512p1[265] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b101010001001,
13'b101010001010,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110101,
13'b1000011110110,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1011011000110,
13'b1011011010101,
13'b1011011010110,
13'b1011011100101,
13'b1011011100110,
13'b1011011110101,
13'b1011011110110,
13'b1100011010101,
13'b1100011010110,
13'b1100011100101,
13'b1100011100110,
13'b1100011110101,
13'b1100011110110,
13'b1101011100101,
13'b1101011110101: edge_mask_reg_512p1[266] <= 1'b1;
 		default: edge_mask_reg_512p1[266] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111011,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101010,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110110,
13'b1001010110110,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1100011010101,
13'b1100011010110,
13'b1100011100101,
13'b1100011100110,
13'b1100011110101,
13'b1100011110110,
13'b1101011010110,
13'b1101011100101,
13'b1101011100110,
13'b1101011110101,
13'b1101011110110: edge_mask_reg_512p1[267] <= 1'b1;
 		default: edge_mask_reg_512p1[267] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101010,
13'b11100101011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b110010001010,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1001010110101,
13'b1001010110110,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1010010110110,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011110101,
13'b1100011110110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100101,
13'b1101011100110,
13'b1101011110101,
13'b1101011110110: edge_mask_reg_512p1[268] <= 1'b1;
 		default: edge_mask_reg_512p1[268] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101010,
13'b11100101011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011110101,
13'b1100011110110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100101,
13'b1101011100110,
13'b1101011110101,
13'b1101011110110,
13'b1110011100110: edge_mask_reg_512p1[269] <= 1'b1;
 		default: edge_mask_reg_512p1[269] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101010,
13'b11100101011,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101010,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101010,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001010,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100101,
13'b1101011100110,
13'b1101011110110,
13'b1110011010110,
13'b1110011100110: edge_mask_reg_512p1[270] <= 1'b1;
 		default: edge_mask_reg_512p1[270] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111011,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101011,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101010,
13'b101001111010,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100001010,
13'b1000010100111,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001010,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011010,
13'b1000011100111,
13'b1000011101000,
13'b1001010100110,
13'b1001010100111,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1010010100110,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110110,
13'b1101011000110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100101,
13'b1101011100110,
13'b1101011110110,
13'b1110011010110,
13'b1110011100110: edge_mask_reg_512p1[271] <= 1'b1;
 		default: edge_mask_reg_512p1[271] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111011,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100001010,
13'b1000010100110,
13'b1000010100111,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011010,
13'b1000011100111,
13'b1000011101000,
13'b1001010100110,
13'b1001010100111,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100111,
13'b1001011101000,
13'b1010010100110,
13'b1010010100111,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100110,
13'b1010011100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1100010110110,
13'b1100010110111,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110110,
13'b1101011000110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100110,
13'b1101011110110,
13'b1110011010110,
13'b1110011100110: edge_mask_reg_512p1[272] <= 1'b1;
 		default: edge_mask_reg_512p1[272] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011010,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011011010,
13'b1000011100111,
13'b1000011101000,
13'b1001010100110,
13'b1001010100111,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100111,
13'b1001011101000,
13'b1010010100110,
13'b1010010100111,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100111,
13'b1011010100110,
13'b1011010100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100110,
13'b1011011100111,
13'b1100010110110,
13'b1100010110111,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1101011000110,
13'b1101011000111,
13'b1101011010110,
13'b1101011010111,
13'b1101011100110,
13'b1110011000110,
13'b1110011010110,
13'b1110011100110: edge_mask_reg_512p1[273] <= 1'b1;
 		default: edge_mask_reg_512p1[273] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101011,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011010,
13'b11100011011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b110001111010,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011010,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101000,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b1000010100111,
13'b1000010101000,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011011010,
13'b1000011101000,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100111,
13'b1001011101000,
13'b1010010100110,
13'b1010010100111,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100111,
13'b1011010100110,
13'b1011010100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100110,
13'b1011011100111,
13'b1100010110110,
13'b1100010110111,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100110,
13'b1101010110110,
13'b1101011000110,
13'b1101011000111,
13'b1101011010110,
13'b1101011010111,
13'b1101011100110,
13'b1110011000110,
13'b1110011010110,
13'b1110011100110: edge_mask_reg_512p1[274] <= 1'b1;
 		default: edge_mask_reg_512p1[274] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011010,
13'b11100011011,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011010,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b111010001001,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101000,
13'b111011101010,
13'b111011111010,
13'b1000010100111,
13'b1000010101000,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011101000,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010111,
13'b1001011011000,
13'b1001011101000,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1011010100110,
13'b1011010100111,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100110,
13'b1100010100111,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100110,
13'b1101010110110,
13'b1101010110111,
13'b1101011000110,
13'b1101011000111,
13'b1101011010110,
13'b1101011010111,
13'b1101011100110,
13'b1110011000110,
13'b1110011010110,
13'b1110011010111: edge_mask_reg_512p1[275] <= 1'b1;
 		default: edge_mask_reg_512p1[275] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011010,
13'b11100011011,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011010,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011010,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101010,
13'b111011111010,
13'b1000010011000,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1001010011000,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010111,
13'b1001011011000,
13'b1010010010111,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010111,
13'b1010011011000,
13'b1011010010111,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1100010100111,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100110,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010110,
13'b1101011010111,
13'b1101011100110,
13'b1110010110110,
13'b1110011000110,
13'b1110011000111,
13'b1110011010110,
13'b1110011010111: edge_mask_reg_512p1[276] <= 1'b1;
 		default: edge_mask_reg_512p1[276] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111010,
13'b10010111011,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b10100011011,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011011,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011010,
13'b101001101010,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011010,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b111010001010,
13'b111010001011,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101010,
13'b111011101011,
13'b111011111010,
13'b111011111011,
13'b1000010011000,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011011000,
13'b1001010011000,
13'b1001010100111,
13'b1001010101000,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010111,
13'b1001011011000,
13'b1010010010111,
13'b1010010011000,
13'b1010010100111,
13'b1010010101000,
13'b1010010110111,
13'b1010010111000,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010111,
13'b1010011011000,
13'b1011010010111,
13'b1011010100111,
13'b1011010101000,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1100010010111,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1101010100111,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010110,
13'b1101011010111,
13'b1110010110110,
13'b1110010110111,
13'b1110011000110,
13'b1110011000111,
13'b1110011010110,
13'b1110011010111: edge_mask_reg_512p1[277] <= 1'b1;
 		default: edge_mask_reg_512p1[277] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111010,
13'b10010111011,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b10100011011,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011011,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011010,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001010,
13'b110100001011,
13'b111001111010,
13'b111001111011,
13'b111010001010,
13'b111010001011,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101010,
13'b111011101011,
13'b111011111010,
13'b111011111011,
13'b1000010011000,
13'b1000010011001,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011011000,
13'b1001010010111,
13'b1001010011000,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010111,
13'b1001011011000,
13'b1010010010111,
13'b1010010011000,
13'b1010010100111,
13'b1010010101000,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010111,
13'b1010011011000,
13'b1011010010111,
13'b1011010011000,
13'b1011010100111,
13'b1011010101000,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010111,
13'b1011011011000,
13'b1100010010111,
13'b1100010011000,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1101010100111,
13'b1101010101000,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1110010110110,
13'b1110010110111,
13'b1110011000110,
13'b1110011000111,
13'b1110011010110,
13'b1110011010111,
13'b1111010110110,
13'b1111010110111,
13'b1111011000110: edge_mask_reg_512p1[278] <= 1'b1;
 		default: edge_mask_reg_512p1[278] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b10100011011,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b110001101010,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001010,
13'b110100001011,
13'b111001111010,
13'b111001111011,
13'b111010001010,
13'b111010001011,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101010,
13'b111011101011,
13'b111011111010,
13'b1000010011000,
13'b1000010011001,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011001000,
13'b1000011001001,
13'b1000011011000,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011001000,
13'b1001011001001,
13'b1001011011000,
13'b1010010010111,
13'b1010010011000,
13'b1010010100111,
13'b1010010101000,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010111,
13'b1010011011000,
13'b1011010010111,
13'b1011010011000,
13'b1011010100111,
13'b1011010101000,
13'b1011010110111,
13'b1011010111000,
13'b1011011000111,
13'b1011011001000,
13'b1011011010111,
13'b1011011011000,
13'b1100010010111,
13'b1100010011000,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010111,
13'b1100011011000,
13'b1101010010111,
13'b1101010011000,
13'b1101010100111,
13'b1101010101000,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1110010110110,
13'b1110010110111,
13'b1110011000110,
13'b1110011000111,
13'b1111010110110,
13'b1111010110111,
13'b1111011000110,
13'b1111011000111: edge_mask_reg_512p1[279] <= 1'b1;
 		default: edge_mask_reg_512p1[279] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011011,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001010,
13'b100100001011,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001010,
13'b101100001011,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111010,
13'b110011111011,
13'b110100001010,
13'b110100001011,
13'b111001111010,
13'b111001111011,
13'b111010001010,
13'b111010001011,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101010,
13'b111011101011,
13'b1000010011000,
13'b1000010011001,
13'b1000010101000,
13'b1000010101001,
13'b1000010111000,
13'b1000010111001,
13'b1000011001000,
13'b1000011001001,
13'b1000011011000,
13'b1001010011000,
13'b1001010011001,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010111000,
13'b1001010111001,
13'b1001011001000,
13'b1001011001001,
13'b1001011011000,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011011000,
13'b1011010010111,
13'b1011010011000,
13'b1011010100111,
13'b1011010101000,
13'b1011010110111,
13'b1011010111000,
13'b1011011000111,
13'b1011011001000,
13'b1011011010111,
13'b1011011011000,
13'b1100010010111,
13'b1100010011000,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010111,
13'b1100011011000,
13'b1101010010111,
13'b1101010011000,
13'b1101010100110,
13'b1101010100111,
13'b1101010101000,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010111,
13'b1110010100110,
13'b1110010100111,
13'b1110010110110,
13'b1110010110111,
13'b1110011000110,
13'b1110011000111,
13'b1111010110111,
13'b1111011000111: edge_mask_reg_512p1[280] <= 1'b1;
 		default: edge_mask_reg_512p1[280] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011011,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001010,
13'b11100001011,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001010,
13'b100100001011,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001010,
13'b101100001011,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111010,
13'b110011111011,
13'b110100001010,
13'b110100001011,
13'b111001111010,
13'b111001111011,
13'b111010001010,
13'b111010001011,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011011010,
13'b111011011011,
13'b111011101010,
13'b111011101011,
13'b1000010011000,
13'b1000010011001,
13'b1000010101000,
13'b1000010101001,
13'b1000010111000,
13'b1000010111001,
13'b1000011001000,
13'b1000011001001,
13'b1000011011000,
13'b1001010011000,
13'b1001010011001,
13'b1001010101000,
13'b1001010101001,
13'b1001010111000,
13'b1001010111001,
13'b1001011001000,
13'b1001011001001,
13'b1001011011000,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011011000,
13'b1011010010111,
13'b1011010011000,
13'b1011010011001,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010110111,
13'b1011010111000,
13'b1011010111001,
13'b1011011000111,
13'b1011011001000,
13'b1011011001001,
13'b1011011011000,
13'b1100010010111,
13'b1100010011000,
13'b1100010100111,
13'b1100010101000,
13'b1100010110111,
13'b1100010111000,
13'b1100011000111,
13'b1100011001000,
13'b1101010010111,
13'b1101010011000,
13'b1101010100110,
13'b1101010100111,
13'b1101010101000,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1110010100110,
13'b1110010100111,
13'b1110010101000,
13'b1110010110110,
13'b1110010110111,
13'b1110010111000,
13'b1110011000111,
13'b1111010100111,
13'b1111010110111,
13'b1111011000111: edge_mask_reg_512p1[281] <= 1'b1;
 		default: edge_mask_reg_512p1[281] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011010101,
13'b10011010110,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101001001,
13'b110101001010,
13'b111001111010,
13'b111001111011,
13'b111010001010,
13'b111010001011,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000010011000,
13'b1000010011001,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011011010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1001010011000,
13'b1001010011001,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011010010111,
13'b1011010011000,
13'b1011010011001,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011010111001,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011001001,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1100010010111,
13'b1100010011000,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1100100000101,
13'b1101010010111,
13'b1101010011000,
13'b1101010100110,
13'b1101010100111,
13'b1101010101000,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1101011100101,
13'b1101011100110,
13'b1101011110101,
13'b1101011110110,
13'b1110010100110,
13'b1110010100111,
13'b1110010101000,
13'b1110010110110,
13'b1110010110111,
13'b1110010111000,
13'b1110011000110,
13'b1110011000111,
13'b1110011010110,
13'b1110011010111,
13'b1110011100110,
13'b1111010100111,
13'b1111010110110,
13'b1111010110111,
13'b1111011000110,
13'b1111011000111: edge_mask_reg_512p1[282] <= 1'b1;
 		default: edge_mask_reg_512p1[282] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011011,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001010,
13'b11100001011,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001010,
13'b101100001011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111001111011,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010011001,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011010111001,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011001001,
13'b1011011011000,
13'b1100010010101,
13'b1100010010110,
13'b1100010010111,
13'b1100010011000,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1101010010100,
13'b1101010010101,
13'b1101010010110,
13'b1101010010111,
13'b1101010011000,
13'b1101010100100,
13'b1101010100101,
13'b1101010100110,
13'b1101010100111,
13'b1101010101000,
13'b1101010110100,
13'b1101010110101,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000101,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1110010010100,
13'b1110010010101,
13'b1110010100100,
13'b1110010100101,
13'b1110010100110,
13'b1110010100111,
13'b1110010101000,
13'b1110010110100,
13'b1110010110101,
13'b1110010110110,
13'b1110010110111,
13'b1110010111000,
13'b1110011000101,
13'b1110011000110,
13'b1110011000111,
13'b1111010100101,
13'b1111010100110,
13'b1111010100111,
13'b1111010110101,
13'b1111010110110,
13'b1111010110111,
13'b1111011000110,
13'b1111011000111: edge_mask_reg_512p1[283] <= 1'b1;
 		default: edge_mask_reg_512p1[283] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011001,
13'b11101011010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101000101,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1000100100011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011,
13'b1001100100011: edge_mask_reg_512p1[284] <= 1'b1;
 		default: edge_mask_reg_512p1[284] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b101011000100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b111101001010,
13'b1000011100011,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011,
13'b1001100100011: edge_mask_reg_512p1[285] <= 1'b1;
 		default: edge_mask_reg_512p1[285] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101001,
13'b11101101010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010100,
13'b100101010101,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b100101101010,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b110011010100,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101011001,
13'b110101011010,
13'b111011011001,
13'b111011011010,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101001001,
13'b111101001010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011,
13'b1001100100011,
13'b1001100110011: edge_mask_reg_512p1[286] <= 1'b1;
 		default: edge_mask_reg_512p1[286] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100011010,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111001,
13'b100101111010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101011001,
13'b111101011010,
13'b1000011110011,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100: edge_mask_reg_512p1[287] <= 1'b1;
 		default: edge_mask_reg_512p1[287] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100101010,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111001,
13'b100101111010,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100100,
13'b101101100101,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b110011100100,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100100,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101011010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101000100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1010100010011,
13'b1010100110011: edge_mask_reg_512p1[288] <= 1'b1;
 		default: edge_mask_reg_512p1[288] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001010,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001001,
13'b100110001010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100100,
13'b110101100101,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101101001,
13'b111101101010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100: edge_mask_reg_512p1[289] <= 1'b1;
 		default: edge_mask_reg_512p1[289] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100111010,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100101,
13'b11101100110,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001001,
13'b100110001010,
13'b101011101001,
13'b101011101010,
13'b101011110101,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101101001,
13'b111101101010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100: edge_mask_reg_512p1[290] <= 1'b1;
 		default: edge_mask_reg_512p1[290] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000101,
13'b100100000110,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011001,
13'b100110011010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101111001,
13'b111101111010,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100101,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100: edge_mask_reg_512p1[291] <= 1'b1;
 		default: edge_mask_reg_512p1[291] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1101001010,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011001,
13'b100110011010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101111001,
13'b111101111010,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110100,
13'b1000101110101,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100: edge_mask_reg_512p1[292] <= 1'b1;
 		default: edge_mask_reg_512p1[292] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000100,
13'b110110000101,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110001001,
13'b111110001010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110100,
13'b1000101110101,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100: edge_mask_reg_512p1[293] <= 1'b1;
 		default: edge_mask_reg_512p1[293] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b111110011010,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000110000101,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1010101000100,
13'b1010101010100,
13'b1010101100100,
13'b1010101110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100: edge_mask_reg_512p1[294] <= 1'b1;
 		default: edge_mask_reg_512p1[294] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110100011001,
13'b110100011010,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110011001,
13'b111110011010,
13'b1000100110101,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000101,
13'b1000110000110,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1010101000100,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101110100,
13'b1010101110101,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[295] <= 1'b1;
 		default: edge_mask_reg_512p1[295] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b111110101010,
13'b1000100110101,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010101,
13'b1000110010110,
13'b1001101000101,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110010101,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010110000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[296] <= 1'b1;
 		default: edge_mask_reg_512p1[296] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b101111001001,
13'b101111001010,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100101,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110101001,
13'b111110101010,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010101,
13'b1000110010110,
13'b1001101000101,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010101,
13'b1001110010110,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010110000100,
13'b1010110000101,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100,
13'b1011110000100: edge_mask_reg_512p1[297] <= 1'b1;
 		default: edge_mask_reg_512p1[297] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001001,
13'b101111001010,
13'b110100111001,
13'b110100111010,
13'b110101000110,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100101,
13'b110110100110,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b110111001001,
13'b110111001010,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110100110,
13'b111110101001,
13'b111110101010,
13'b111110111001,
13'b111110111010,
13'b1000101000101,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100101,
13'b1000110100110,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100101,
13'b1001110100110,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010110000100,
13'b1010110000101,
13'b1010110010100,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101: edge_mask_reg_512p1[298] <= 1'b1;
 		default: edge_mask_reg_512p1[298] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001001,
13'b10110001010,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001001,
13'b101111001010,
13'b101111011001,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b110111001001,
13'b110111001010,
13'b111101001001,
13'b111101001010,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101001,
13'b111110101010,
13'b111110111001,
13'b111110111010,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100101,
13'b1000110100110,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100101,
13'b1001110100110,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010110000100,
13'b1010110000101,
13'b1010110010100,
13'b1010110010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1011110010100,
13'b1011110010101,
13'b1100101110100,
13'b1100110010100: edge_mask_reg_512p1[299] <= 1'b1;
 		default: edge_mask_reg_512p1[299] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001001,
13'b10110001010,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011001,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111001001,
13'b110111001010,
13'b110111011001,
13'b110111011010,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101001,
13'b111110101010,
13'b111110110101,
13'b111110110110,
13'b111110111001,
13'b111110111010,
13'b111111001001,
13'b111111001010,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110101,
13'b1001110110110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1011110010100,
13'b1011110010101,
13'b1011110100100,
13'b1100101110100,
13'b1100101110101,
13'b1100110000100,
13'b1100110000101,
13'b1100110010100,
13'b1100110010101: edge_mask_reg_512p1[300] <= 1'b1;
 		default: edge_mask_reg_512p1[300] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001010,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10110001001,
13'b10110001010,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011001,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b110101100110,
13'b110101100111,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111001001,
13'b110111001010,
13'b110111011001,
13'b110111011010,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111001,
13'b111110111010,
13'b111111001001,
13'b111111001010,
13'b1000101100101,
13'b1000101100110,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110101,
13'b1001110110110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110101,
13'b1010110110110,
13'b1011101110100,
13'b1011110000100,
13'b1011110000101,
13'b1011110010100,
13'b1011110010101,
13'b1011110100100,
13'b1011110100101,
13'b1100110000100,
13'b1100110000101,
13'b1100110010100,
13'b1100110010101,
13'b1100110100100,
13'b1100110100101: edge_mask_reg_512p1[301] <= 1'b1;
 		default: edge_mask_reg_512p1[301] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001001,
13'b10110001010,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111011001,
13'b110111011010,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000101,
13'b111111000110,
13'b111111001001,
13'b111111001010,
13'b111111011001,
13'b111111011010,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000101,
13'b1000111000110,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000101,
13'b1001111000110,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000101,
13'b1010111000110,
13'b1011110000100,
13'b1011110000101,
13'b1011110010100,
13'b1011110010101,
13'b1011110100100,
13'b1011110100101,
13'b1011110110100,
13'b1011110110101,
13'b1100110000100,
13'b1100110000101,
13'b1100110010100,
13'b1100110010101,
13'b1100110100100,
13'b1100110100101: edge_mask_reg_512p1[302] <= 1'b1;
 		default: edge_mask_reg_512p1[302] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b110101110110,
13'b110101110111,
13'b110101111001,
13'b110101111010,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111011001,
13'b110111011010,
13'b111101101001,
13'b111101101010,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111011001,
13'b111111011010,
13'b1000101110101,
13'b1000101110110,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000101,
13'b1001111000110,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000101,
13'b1010111000110,
13'b1011110010100,
13'b1011110010101,
13'b1011110100100,
13'b1011110100101,
13'b1011110110100,
13'b1011110110101,
13'b1100110010101,
13'b1100110100101,
13'b1100110110101: edge_mask_reg_512p1[303] <= 1'b1;
 		default: edge_mask_reg_512p1[303] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011001,
13'b110111011010,
13'b111101111001,
13'b111101111010,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011001,
13'b111111011010,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1001110000101,
13'b1001110000110,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100101,
13'b1001110100110,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010101,
13'b1001111010110,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010101,
13'b1010111010110,
13'b1011110010100,
13'b1011110010101,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011111000100,
13'b1011111000101,
13'b1100110010101,
13'b1100110100101,
13'b1100110110101,
13'b1100111000101: edge_mask_reg_512p1[304] <= 1'b1;
 		default: edge_mask_reg_512p1[304] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101111001,
13'b111101111010,
13'b111110000110,
13'b111110001001,
13'b111110001010,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b1000110000101,
13'b1000110000110,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1001110000101,
13'b1001110000110,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110101,
13'b1001110110110,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1010110010101,
13'b1010110010110,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010101,
13'b1010111010110,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1100110100101,
13'b1100110110101,
13'b1100111000101: edge_mask_reg_512p1[305] <= 1'b1;
 		default: edge_mask_reg_512p1[305] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110001001,
13'b111110001010,
13'b111110010110,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b1000110010110,
13'b1000110010111,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100110,
13'b1000111100111,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100110,
13'b1010110010110,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100110,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111010101,
13'b1011111010110,
13'b1100110100101,
13'b1100110110101,
13'b1100111000101,
13'b1100111010101,
13'b1101110100101,
13'b1101110110101,
13'b1101111000101: edge_mask_reg_512p1[306] <= 1'b1;
 		default: edge_mask_reg_512p1[306] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b111110011010,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b1000110010110,
13'b1000110010111,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110100110,
13'b1001110100111,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100110,
13'b1001111100111,
13'b1010110100110,
13'b1010110100111,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100110,
13'b1010111100111,
13'b1011110100110,
13'b1011110110101,
13'b1011110110110,
13'b1011111000101,
13'b1011111000110,
13'b1011111010101,
13'b1011111010110,
13'b1011111100110,
13'b1100110110101,
13'b1100110110110,
13'b1100111000101,
13'b1100111000110,
13'b1100111010101,
13'b1100111010110,
13'b1101110110101,
13'b1101111000101,
13'b1101111010101: edge_mask_reg_512p1[307] <= 1'b1;
 		default: edge_mask_reg_512p1[307] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110011001,
13'b111110011010,
13'b111110100110,
13'b111110100111,
13'b111110101001,
13'b111110101010,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b1000110100110,
13'b1000110100111,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110100110,
13'b1001110100111,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100110,
13'b1001111100111,
13'b1010110100110,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1011110100110,
13'b1011110110101,
13'b1011110110110,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1100110110101,
13'b1100110110110,
13'b1100111000101,
13'b1100111000110,
13'b1100111010101,
13'b1100111010110,
13'b1100111100101,
13'b1100111100110,
13'b1101110110101,
13'b1101111000101,
13'b1101111010101,
13'b1101111100101: edge_mask_reg_512p1[308] <= 1'b1;
 		default: edge_mask_reg_512p1[308] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101101000,
13'b101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b111110101010,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000110100111,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110110110,
13'b1001110110111,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100110,
13'b1001111100111,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1011110110110,
13'b1011110110111,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1011111110111,
13'b1100111000101,
13'b1100111000110,
13'b1100111010101,
13'b1100111010110,
13'b1100111100101,
13'b1100111100110,
13'b1101111000101,
13'b1101111010101,
13'b1101111100101: edge_mask_reg_512p1[309] <= 1'b1;
 		default: edge_mask_reg_512p1[309] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101101001,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110101001,
13'b111110101010,
13'b111110110110,
13'b111110110111,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000110110110,
13'b1000110110111,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110110110,
13'b1001110110111,
13'b1001111000110,
13'b1001111000111,
13'b1001111010110,
13'b1001111010111,
13'b1001111100110,
13'b1001111100111,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110111,
13'b1011110110110,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1011111110111,
13'b1100111000101,
13'b1100111000110,
13'b1100111010101,
13'b1100111010110,
13'b1100111100101,
13'b1100111100110,
13'b1100111110101,
13'b1100111110110,
13'b1101111000101,
13'b1101111010101,
13'b1101111010110,
13'b1101111100101,
13'b1101111100110,
13'b1101111110101,
13'b1101111110110: edge_mask_reg_512p1[310] <= 1'b1;
 		default: edge_mask_reg_512p1[310] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110101001,
13'b111110101010,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001111000110,
13'b1001111000111,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110111,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1011111110111,
13'b1100111010101,
13'b1100111010110,
13'b1100111010111,
13'b1100111100101,
13'b1100111100110,
13'b1100111100111,
13'b1100111110101,
13'b1100111110110,
13'b1100111110111,
13'b1101111010101,
13'b1101111010110,
13'b1101111100101,
13'b1101111100110,
13'b1101111110101,
13'b1101111110110: edge_mask_reg_512p1[311] <= 1'b1;
 		default: edge_mask_reg_512p1[311] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1110001001,
13'b1110001010,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110111001,
13'b111110111010,
13'b111111000111,
13'b111111001001,
13'b111111001010,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000111000111,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001111000110,
13'b1001111000111,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1011111110111,
13'b1100111010101,
13'b1100111010110,
13'b1100111010111,
13'b1100111100101,
13'b1100111100110,
13'b1100111100111,
13'b1100111110101,
13'b1100111110110,
13'b1100111110111,
13'b1101111010101,
13'b1101111100101,
13'b1101111100110,
13'b1101111110101,
13'b1101111110110: edge_mask_reg_512p1[312] <= 1'b1;
 		default: edge_mask_reg_512p1[312] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110011010,
13'b10110101001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110111001,
13'b111110111010,
13'b111111001001,
13'b111111001010,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010111010110,
13'b1010111010111,
13'b1010111100110,
13'b1010111100111,
13'b1010111110111,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1011111110111,
13'b1100111010110,
13'b1100111010111,
13'b1100111100101,
13'b1100111100110,
13'b1100111100111,
13'b1100111110101,
13'b1100111110110,
13'b1100111110111,
13'b1101111100101,
13'b1101111100110,
13'b1101111110101,
13'b1101111110110,
13'b1110111100110,
13'b1110111110110: edge_mask_reg_512p1[313] <= 1'b1;
 		default: edge_mask_reg_512p1[313] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110011010,
13'b10110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111111001001,
13'b111111001010,
13'b111111010111,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000111100111,
13'b1000111101000,
13'b1001111010110,
13'b1001111010111,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010111010110,
13'b1010111010111,
13'b1010111100110,
13'b1010111100111,
13'b1010111101000,
13'b1010111110111,
13'b1010111111000,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1011111110111,
13'b1100111100110,
13'b1100111100111,
13'b1100111110101,
13'b1100111110110,
13'b1100111110111,
13'b1101111110101,
13'b1101111110110,
13'b1110111110110: edge_mask_reg_512p1[314] <= 1'b1;
 		default: edge_mask_reg_512p1[314] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101010101001,
13'b101010110100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111011001001,
13'b111011001010,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000011010011,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001011100011,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110111,
13'b1010111111000,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1011110010100,
13'b1011110010101,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1011111110111,
13'b1100101110100,
13'b1100101110101,
13'b1100110000100,
13'b1100110000101,
13'b1100110010100,
13'b1100110010101,
13'b1100110100100,
13'b1100110100101,
13'b1100110110101,
13'b1100110110110,
13'b1100111000101,
13'b1100111000110,
13'b1100111010101,
13'b1100111010110,
13'b1100111010111,
13'b1100111100101,
13'b1100111100110,
13'b1100111100111,
13'b1100111110101,
13'b1100111110110,
13'b1100111110111,
13'b1101110100101,
13'b1101110110101,
13'b1101111000101,
13'b1101111010101,
13'b1101111010110,
13'b1101111100101,
13'b1101111100110,
13'b1101111110101,
13'b1101111110110,
13'b1110111100110,
13'b1110111110110: edge_mask_reg_512p1[315] <= 1'b1;
 		default: edge_mask_reg_512p1[315] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111111001010,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110111,
13'b1010111111000,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1011111110111,
13'b1100111100110,
13'b1100111100111,
13'b1100111110101,
13'b1100111110110,
13'b1100111110111,
13'b1101111110101,
13'b1101111110110,
13'b1110111110101,
13'b1110111110110: edge_mask_reg_512p1[316] <= 1'b1;
 		default: edge_mask_reg_512p1[316] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010110100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b1000011010011,
13'b1000011100011,
13'b1000011110011,
13'b1000100000011,
13'b1000100010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100010011: edge_mask_reg_512p1[317] <= 1'b1;
 		default: edge_mask_reg_512p1[317] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011111010,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001001,
13'b11101001010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100111001,
13'b110100111010,
13'b111010111001,
13'b111010111010,
13'b111011001001,
13'b111011001010,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1001011010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011: edge_mask_reg_512p1[318] <= 1'b1;
 		default: edge_mask_reg_512p1[318] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011101010,
13'b1011111001,
13'b1011111010,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110110,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b100010011001,
13'b100010011010,
13'b100010100100,
13'b100010100101,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b111010110100,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b1000011000011,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1001011000011,
13'b1001011010011,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011: edge_mask_reg_512p1[319] <= 1'b1;
 		default: edge_mask_reg_512p1[319] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011101010,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110110,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100101,
13'b11010100110,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111001,
13'b11100111010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100100,
13'b100010100101,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b1000011000011,
13'b1000011000100,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100: edge_mask_reg_512p1[320] <= 1'b1;
 		default: edge_mask_reg_512p1[320] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011011010,
13'b1011101001,
13'b1011101010,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010100,
13'b100100010101,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101001,
13'b100100101010,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010100100,
13'b111010100101,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b1000010110011,
13'b1000010110100,
13'b1000011000011,
13'b1000011000100,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1001010110011,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1010011000011,
13'b1010011100011: edge_mask_reg_512p1[321] <= 1'b1;
 		default: edge_mask_reg_512p1[321] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011011010,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101001,
13'b100100101010,
13'b101010001001,
13'b101010001010,
13'b101010010100,
13'b101010010101,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b111010010100,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b1000010110011,
13'b1000010110100,
13'b1000011000011,
13'b1000011000100,
13'b1000011010011,
13'b1000011010100,
13'b1000011100011,
13'b1000011100100,
13'b1001010110011,
13'b1001010110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100: edge_mask_reg_512p1[322] <= 1'b1;
 		default: edge_mask_reg_512p1[322] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1011001010,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011001,
13'b100100011010,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b111010001001,
13'b111010010100,
13'b111010010101,
13'b111010011001,
13'b111010011010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1001010100011,
13'b1001010100100,
13'b1001010110011,
13'b1001010110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100: edge_mask_reg_512p1[323] <= 1'b1;
 		default: edge_mask_reg_512p1[323] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1011001010,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011001,
13'b100100011010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b110001111001,
13'b110001111010,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b111010000100,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100101,
13'b1001010100011,
13'b1001010100100,
13'b1001010110011,
13'b1001010110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100: edge_mask_reg_512p1[324] <= 1'b1;
 		default: edge_mask_reg_512p1[324] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010111010,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000101,
13'b100010000110,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001001,
13'b100100001010,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b1000010000101,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1001010010011,
13'b1001010010100,
13'b1001010100011,
13'b1001010100100,
13'b1001010110011,
13'b1001010110100,
13'b1001011000011,
13'b1001011000100,
13'b1001011010011,
13'b1001011010100,
13'b1010010010011,
13'b1010010010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100: edge_mask_reg_512p1[325] <= 1'b1;
 		default: edge_mask_reg_512p1[325] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001010,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001001,
13'b100100001010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b110001101001,
13'b110001101010,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001110100,
13'b111001110101,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011101001,
13'b111011101010,
13'b1000010000100,
13'b1000010000101,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010100,
13'b1000011010101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1010010010011,
13'b1010010010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100: edge_mask_reg_512p1[326] <= 1'b1;
 		default: edge_mask_reg_512p1[326] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110101,
13'b101001110110,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b1000001110101,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010100,
13'b1000011010101,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1010010000100,
13'b1010010010100,
13'b1010010100100,
13'b1010010110100,
13'b1011010010100,
13'b1011010100100,
13'b1011010110100: edge_mask_reg_512p1[327] <= 1'b1;
 		default: edge_mask_reg_512p1[327] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111010,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b101011111010,
13'b110001011001,
13'b110001011010,
13'b110001100101,
13'b110001100110,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001100101,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010100100,
13'b1010010100101,
13'b1010010110100,
13'b1011010000100,
13'b1011010010100,
13'b1011010100100,
13'b1011010110100: edge_mask_reg_512p1[328] <= 1'b1;
 		default: edge_mask_reg_512p1[328] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001010,
13'b1001111001,
13'b1010001010,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b10001101000,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101001,
13'b100011101010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100101,
13'b101001100110,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b110001001010,
13'b110001011001,
13'b110001011010,
13'b110001100101,
13'b110001100110,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1001001100101,
13'b1001001110100,
13'b1001001110101,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110101,
13'b1010001110100,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1010010100100,
13'b1010010100101,
13'b1011010000100,
13'b1011010010100,
13'b1011010100100: edge_mask_reg_512p1[329] <= 1'b1;
 		default: edge_mask_reg_512p1[329] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b1001111001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b10001101000,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101001,
13'b100011101010,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011001,
13'b101011011010,
13'b110001001001,
13'b110001001010,
13'b110001010110,
13'b110001011001,
13'b110001011010,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001001,
13'b110011001010,
13'b110011011001,
13'b110011011010,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011001001,
13'b111011001010,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110101,
13'b1000010110110,
13'b1001001100101,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110101,
13'b1010001110100,
13'b1010001110101,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1010010100100,
13'b1010010100101,
13'b1011001110100,
13'b1011010000100,
13'b1011010010100,
13'b1011010100100: edge_mask_reg_512p1[330] <= 1'b1;
 		default: edge_mask_reg_512p1[330] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111010,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011001,
13'b101011011010,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b110001010101,
13'b110001010110,
13'b110001011001,
13'b110001011010,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100101,
13'b1000010100110,
13'b1000010110101,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100101,
13'b1001010100110,
13'b1010001100100,
13'b1010001100101,
13'b1010001110100,
13'b1010001110101,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1011001100100,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101: edge_mask_reg_512p1[331] <= 1'b1;
 		default: edge_mask_reg_512p1[331] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001001,
13'b101011001010,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b111001000110,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100101,
13'b1000010100110,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100101,
13'b1001010100110,
13'b1010001100100,
13'b1010001100101,
13'b1010001110100,
13'b1010001110101,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1011001100100,
13'b1011001100101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1100001100100,
13'b1100010000100: edge_mask_reg_512p1[332] <= 1'b1;
 		default: edge_mask_reg_512p1[332] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101011001001,
13'b101011001010,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001001,
13'b110001001010,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010101001,
13'b111010101010,
13'b1000001000101,
13'b1000001000110,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010101,
13'b1000010010110,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010101,
13'b1001010010110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001100100,
13'b1011001100101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1100001100100,
13'b1100001100101,
13'b1100001110100,
13'b1100001110101,
13'b1100010000100: edge_mask_reg_512p1[333] <= 1'b1;
 		default: edge_mask_reg_512p1[333] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001010,
13'b10011001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010110,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b111000110110,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010101,
13'b1000010010110,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010101,
13'b1001010010110,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001100100,
13'b1011001100101,
13'b1011001110100,
13'b1011001110101,
13'b1100001010100,
13'b1100001010101,
13'b1100001100100,
13'b1100001100101,
13'b1100001110100,
13'b1100001110101: edge_mask_reg_512p1[334] <= 1'b1;
 		default: edge_mask_reg_512p1[334] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b110000110110,
13'b110000110111,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b1000000110101,
13'b1000000110110,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1001000110101,
13'b1001000110110,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000101,
13'b1001010000110,
13'b1010000110101,
13'b1010000110110,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000101,
13'b1010010000110,
13'b1011001000100,
13'b1011001000101,
13'b1011001010100,
13'b1011001010101,
13'b1011001100100,
13'b1011001100101,
13'b1011001110100,
13'b1011001110101,
13'b1100001000101,
13'b1100001010100,
13'b1100001010101,
13'b1100001100100,
13'b1100001100101,
13'b1100001110100,
13'b1100001110101: edge_mask_reg_512p1[335] <= 1'b1;
 		default: edge_mask_reg_512p1[335] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111010,
13'b10010111011,
13'b11001011000,
13'b11001011001,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000110,
13'b110010000111,
13'b110010001001,
13'b110010001010,
13'b110010011001,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b1000000100110,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1001000110101,
13'b1001000110110,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110101,
13'b1001001110110,
13'b1001010000101,
13'b1001010000110,
13'b1010000110101,
13'b1010000110110,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110101,
13'b1010001110110,
13'b1011001000100,
13'b1011001000101,
13'b1011001010100,
13'b1011001010101,
13'b1011001100100,
13'b1011001100101,
13'b1100001000101,
13'b1100001010101,
13'b1100001100101: edge_mask_reg_512p1[336] <= 1'b1;
 		default: edge_mask_reg_512p1[336] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b11001011000,
13'b11001011001,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101010,
13'b11010101011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010011001,
13'b110010011010,
13'b111000100111,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010001001,
13'b111010001010,
13'b1000000100110,
13'b1000000100111,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1001000100101,
13'b1001000100110,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110101,
13'b1001001110110,
13'b1010000100101,
13'b1010000100110,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110101,
13'b1010001110110,
13'b1011000110100,
13'b1011000110101,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100100,
13'b1011001100101,
13'b1100000110101,
13'b1100001000101,
13'b1100001010101,
13'b1100001100101: edge_mask_reg_512p1[337] <= 1'b1;
 		default: edge_mask_reg_512p1[337] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111001,
13'b10111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b11001011000,
13'b11001011001,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110010001001,
13'b110010001010,
13'b110010011001,
13'b110010011010,
13'b111000100111,
13'b111000101000,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001111001,
13'b111001111010,
13'b111010001001,
13'b111010001010,
13'b1000000100110,
13'b1000000100111,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000101,
13'b1001001000110,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110101,
13'b1010000100101,
13'b1010000100110,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100101,
13'b1010001100110,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1100000110101,
13'b1100001000101,
13'b1100001010101: edge_mask_reg_512p1[338] <= 1'b1;
 		default: edge_mask_reg_512p1[338] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b11001011000,
13'b11001011001,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011010,
13'b11010011011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110010001001,
13'b110010001010,
13'b111000100111,
13'b111000101000,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001111001,
13'b111001111010,
13'b1000000100110,
13'b1000000100111,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100110,
13'b1000001100111,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100101,
13'b1001001100110,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001010101,
13'b1010001010110,
13'b1010001100101,
13'b1010001100110,
13'b1011000100101,
13'b1011000100110,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1100000100101,
13'b1100000110101,
13'b1100001000101,
13'b1100001010101,
13'b1101000100101,
13'b1101000110101,
13'b1101001000101,
13'b1101001010101: edge_mask_reg_512p1[339] <= 1'b1;
 		default: edge_mask_reg_512p1[339] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011010,
13'b10010011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110010001001,
13'b110010001010,
13'b111000100111,
13'b111000101000,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001101001,
13'b111001101010,
13'b111001111010,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1000001010110,
13'b1000001010111,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010110,
13'b1001001010111,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001010110,
13'b1010001010111,
13'b1011000010110,
13'b1011000100101,
13'b1011000100110,
13'b1011000110101,
13'b1011000110110,
13'b1011001000101,
13'b1011001000110,
13'b1011001010110,
13'b1100000100101,
13'b1100000100110,
13'b1100000110101,
13'b1100000110110,
13'b1100001000101,
13'b1100001000110,
13'b1101000100101,
13'b1101000110101,
13'b1101001000101: edge_mask_reg_512p1[340] <= 1'b1;
 		default: edge_mask_reg_512p1[340] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001111000,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011010,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001010,
13'b11010001011,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001101001,
13'b111001101010,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1000001010110,
13'b1000001010111,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010110,
13'b1001001010111,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001010110,
13'b1010001010111,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1011001000101,
13'b1011001000110,
13'b1011001010110,
13'b1100000010101,
13'b1100000010110,
13'b1100000100101,
13'b1100000100110,
13'b1100000110101,
13'b1100000110110,
13'b1100001000101,
13'b1100001000110,
13'b1101000010101,
13'b1101000100101,
13'b1101000110101,
13'b1101001000101: edge_mask_reg_512p1[341] <= 1'b1;
 		default: edge_mask_reg_512p1[341] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001010,
13'b10010001011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b100001001000,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001011001,
13'b111001011010,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000110,
13'b1001001000111,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000110,
13'b1010001000111,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1011001000110,
13'b1011001000111,
13'b1100000010101,
13'b1100000010110,
13'b1100000100101,
13'b1100000100110,
13'b1100000110101,
13'b1100000110110,
13'b1101000010101,
13'b1101000100101,
13'b1101000110101: edge_mask_reg_512p1[342] <= 1'b1;
 		default: edge_mask_reg_512p1[342] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001111001,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111010,
13'b11001111011,
13'b100001001000,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111010,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000111,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001011001,
13'b111001011010,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000001000111,
13'b1001000100110,
13'b1001000100111,
13'b1001000110110,
13'b1001000110111,
13'b1001001000110,
13'b1001001000111,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000110,
13'b1010001000111,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1011001000110,
13'b1100000010101,
13'b1100000010110,
13'b1100000100101,
13'b1100000100110,
13'b1100000110101,
13'b1101000010101,
13'b1101000010110,
13'b1101000100101,
13'b1101000100110: edge_mask_reg_512p1[343] <= 1'b1;
 		default: edge_mask_reg_512p1[343] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10001101001,
13'b10001111010,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b101000111000,
13'b101000111001,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101010,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001001001,
13'b111001001010,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110110,
13'b1001000110111,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110110,
13'b1010000110111,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110110,
13'b1011000110111,
13'b1100000010101,
13'b1100000010110,
13'b1100000010111,
13'b1100000100101,
13'b1100000100110,
13'b1100000100111,
13'b1101000010101,
13'b1101000010110,
13'b1101000100101,
13'b1101000100110: edge_mask_reg_512p1[344] <= 1'b1;
 		default: edge_mask_reg_512p1[344] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10001101001,
13'b11001011001,
13'b11001011010,
13'b11001101010,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b101000111001,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101010,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011001,
13'b110001011010,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000111001,
13'b111000111010,
13'b111001001001,
13'b111001001010,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000110111,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110110,
13'b1001000110111,
13'b1010000010111,
13'b1010000100110,
13'b1010000100111,
13'b1010000110110,
13'b1010000110111,
13'b1011000010110,
13'b1011000010111,
13'b1011000100110,
13'b1011000100111,
13'b1100000010101,
13'b1100000010110,
13'b1100000010111,
13'b1100000100110,
13'b1100000100111,
13'b1101000010101,
13'b1101000010110: edge_mask_reg_512p1[345] <= 1'b1;
 		default: edge_mask_reg_512p1[345] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001011001,
13'b11001011010,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b101000111001,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011010,
13'b111000100111,
13'b111000101000,
13'b111000111001,
13'b111000111010,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1010000010111,
13'b1010000100110,
13'b1010000100111,
13'b1011000010110,
13'b1011000010111,
13'b1011000100110,
13'b1011000100111,
13'b1100000010101,
13'b1100000010110,
13'b1100000010111,
13'b1100000100110,
13'b1100000100111,
13'b1101000010101,
13'b1101000010110,
13'b1110000010110: edge_mask_reg_512p1[346] <= 1'b1;
 		default: edge_mask_reg_512p1[346] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001001001,
13'b100001011010,
13'b101000111001,
13'b101001001001,
13'b101001001010,
13'b101001011010,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b111000111001,
13'b111000111010,
13'b1010000010111,
13'b1011000010110,
13'b1011000010111,
13'b1100000010110,
13'b1100000010111: edge_mask_reg_512p1[347] <= 1'b1;
 		default: edge_mask_reg_512p1[347] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111000111011,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001001011,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001011011,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001101011,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111001111011,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000000100111,
13'b1000000101000,
13'b1000000110111,
13'b1000000111000,
13'b1000001000111,
13'b1000001001000,
13'b1000001010111,
13'b1000001011000,
13'b1000001100111,
13'b1000001101000,
13'b1000001110111,
13'b1000001111000,
13'b1000010000111,
13'b1000010001000,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110110,
13'b1001000110111,
13'b1001000111000,
13'b1001001000110,
13'b1001001000111,
13'b1001001001000,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000111,
13'b1001011001000,
13'b1001011010111,
13'b1001011011000,
13'b1001011100111,
13'b1001011101000,
13'b1001011110111,
13'b1001011111000,
13'b1001100000111,
13'b1001100001000,
13'b1001100010111,
13'b1001100011000,
13'b1010000010111,
13'b1010000011000,
13'b1010000100110,
13'b1010000100111,
13'b1010000101000,
13'b1010000110110,
13'b1010000110111,
13'b1010000111000,
13'b1010001000110,
13'b1010001000111,
13'b1010001001000,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1010001100110,
13'b1010001100111,
13'b1010001101000,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010111,
13'b1010100011000,
13'b1011000010110,
13'b1011000010111,
13'b1011000100110,
13'b1011000100111,
13'b1011000110110,
13'b1011000110111,
13'b1011001000110,
13'b1011001000111,
13'b1011001010110,
13'b1011001010111,
13'b1011001100110,
13'b1011001100111,
13'b1011001110110,
13'b1011001110111,
13'b1011010000110,
13'b1011010000111,
13'b1011010010110,
13'b1011010010111,
13'b1011010100110,
13'b1011010100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011010110,
13'b1011011010111,
13'b1011011100110,
13'b1011011100111,
13'b1011011110110,
13'b1011011110111,
13'b1011100000110,
13'b1011100000111,
13'b1011100010110,
13'b1011100010111,
13'b1100000010101,
13'b1100000010110,
13'b1100000010111,
13'b1100000100101,
13'b1100000100110,
13'b1100000100111,
13'b1100000110101,
13'b1100000110110,
13'b1100000110111,
13'b1100001000101,
13'b1100001000110,
13'b1100001000111,
13'b1100001010101,
13'b1100001010110,
13'b1100001010111,
13'b1100001100101,
13'b1100001100110,
13'b1100001100111,
13'b1100001110101,
13'b1100001110110,
13'b1100001110111,
13'b1100010000101,
13'b1100010000110,
13'b1100010000111,
13'b1100010010101,
13'b1100010010110,
13'b1100010010111,
13'b1100010100101,
13'b1100010100110,
13'b1100010100111,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000110,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1101000010101,
13'b1101000010110,
13'b1101000100101,
13'b1101000100110,
13'b1101000110101,
13'b1101000110110,
13'b1101001000101,
13'b1101001000110,
13'b1101001010101,
13'b1101001010110,
13'b1101001010111,
13'b1101001100101,
13'b1101001100110,
13'b1101001100111,
13'b1101001110101,
13'b1101001110110,
13'b1101001110111,
13'b1101010000101,
13'b1101010000110,
13'b1101010000111,
13'b1101010010101,
13'b1101010010110,
13'b1101010010111,
13'b1101010100101,
13'b1101010100110,
13'b1101010100111,
13'b1101010110101,
13'b1101010110110,
13'b1101010110111,
13'b1101011000101,
13'b1101011000110,
13'b1101011000111,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011100110,
13'b1101011100111,
13'b1101011110110,
13'b1101011110111,
13'b1101100000110,
13'b1101100000111,
13'b1101100010111,
13'b1110000010110,
13'b1110000100110,
13'b1110000110110,
13'b1110001000110,
13'b1110001010110,
13'b1110001100110,
13'b1110001110110,
13'b1110010000110,
13'b1110010010110,
13'b1110010100110,
13'b1110010110110,
13'b1110011000110,
13'b1110011010110,
13'b1110011100110,
13'b1110011110110,
13'b1110100000110,
13'b1111011110110,
13'b1111100000110: edge_mask_reg_512p1[348] <= 1'b1;
 		default: edge_mask_reg_512p1[348] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001001001,
13'b101000111000,
13'b101000111001,
13'b101001001001,
13'b101001001010,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001001010,
13'b111000101001,
13'b1010000010111,
13'b1011000010110,
13'b1011000010111,
13'b1100000010110,
13'b1100000010111: edge_mask_reg_512p1[349] <= 1'b1;
 		default: edge_mask_reg_512p1[349] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011010,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100111,
13'b1000011101000,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1001011010111,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1010011010111,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010110,
13'b1011100010111,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1101011100110,
13'b1101011100111,
13'b1101011110101,
13'b1101011110110,
13'b1101011110111,
13'b1101100000101,
13'b1101100000110,
13'b1101100000111,
13'b1101100010111,
13'b1110011110110,
13'b1110100000110,
13'b1111100000110: edge_mask_reg_512p1[350] <= 1'b1;
 		default: edge_mask_reg_512p1[350] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101010,
13'b10101101011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101001010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1001011000101,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1010011010100,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1011011100100,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101: edge_mask_reg_512p1[351] <= 1'b1;
 		default: edge_mask_reg_512p1[351] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101010,
13'b10101101011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b101010011001,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101001010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1001011000101,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1010011010100,
13'b1010011010101,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101: edge_mask_reg_512p1[352] <= 1'b1;
 		default: edge_mask_reg_512p1[352] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101010,
13'b10101101011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101001010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110101,
13'b1100100000101: edge_mask_reg_512p1[353] <= 1'b1;
 		default: edge_mask_reg_512p1[353] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101010,
13'b11100101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101010,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101010,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b111010001001,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b1000010100101,
13'b1000010100110,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1001010100101,
13'b1001010100110,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1010010100101,
13'b1010010100110,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011110101,
13'b1100011110110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100101,
13'b1101011100110,
13'b1101011110101,
13'b1101011110110,
13'b1110011100110: edge_mask_reg_512p1[354] <= 1'b1;
 		default: edge_mask_reg_512p1[354] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001010,
13'b111001000110,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010101001,
13'b111010101010,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1100001100100,
13'b1100001100101,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100010000100,
13'b1100010000101,
13'b1100010000110,
13'b1101001110101,
13'b1101010000101: edge_mask_reg_512p1[355] <= 1'b1;
 		default: edge_mask_reg_512p1[355] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001010,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b1000001000101,
13'b1000001000110,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1011001010100,
13'b1011001010101,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1100001100100,
13'b1100001100101,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100010000101,
13'b1100010000110,
13'b1101001110101,
13'b1101010000101: edge_mask_reg_512p1[356] <= 1'b1;
 		default: edge_mask_reg_512p1[356] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001010,
13'b111000110110,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010110,
13'b1010010010111,
13'b1011001010100,
13'b1011001010101,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1100001010100,
13'b1100001010101,
13'b1100001100100,
13'b1100001100101,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100010000101,
13'b1100010000110,
13'b1101001110101,
13'b1101010000101: edge_mask_reg_512p1[357] <= 1'b1;
 		default: edge_mask_reg_512p1[357] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b110000110110,
13'b110000110111,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001010,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b1000000110101,
13'b1000000110110,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1001000110101,
13'b1001000110110,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1010000110101,
13'b1010000110110,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010110,
13'b1010010010111,
13'b1011001000100,
13'b1011001000101,
13'b1011001010100,
13'b1011001010101,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000101,
13'b1011010000110,
13'b1100001000101,
13'b1100001010101,
13'b1100001100101,
13'b1100001110101,
13'b1100001110110,
13'b1100010000101,
13'b1100010000110,
13'b1101001110101,
13'b1101010000101: edge_mask_reg_512p1[358] <= 1'b1;
 		default: edge_mask_reg_512p1[358] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001101100,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001010,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b1000000100110,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1001000110101,
13'b1001000110110,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010110,
13'b1001010010111,
13'b1010000110101,
13'b1010000110110,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010110,
13'b1010010010111,
13'b1011001000100,
13'b1011001000101,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000101,
13'b1011010000110,
13'b1100001000101,
13'b1100001010101,
13'b1100001100101,
13'b1100001110101,
13'b1100001110110,
13'b1100010000101,
13'b1100010000110,
13'b1101001110101,
13'b1101010000101: edge_mask_reg_512p1[359] <= 1'b1;
 		default: edge_mask_reg_512p1[359] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000110,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000101,
13'b1000110000110,
13'b1001100110101,
13'b1001100110110,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1010101000100,
13'b1010101000101,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1100101010100,
13'b1100101100100: edge_mask_reg_512p1[360] <= 1'b1;
 		default: edge_mask_reg_512p1[360] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b111110011010,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1001100110101,
13'b1001100110110,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1010101000100,
13'b1010101000101,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1100101010100,
13'b1100101100100: edge_mask_reg_512p1[361] <= 1'b1;
 		default: edge_mask_reg_512p1[361] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b110011111001,
13'b110011111010,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100000101,
13'b1000100000110,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110101,
13'b1000101110110,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110101,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1011101000101,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101110100,
13'b1100100100100,
13'b1100100110100,
13'b1100100110101,
13'b1100101000100,
13'b1100101000101: edge_mask_reg_512p1[362] <= 1'b1;
 		default: edge_mask_reg_512p1[362] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101010,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110011111001,
13'b110011111010,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100000101,
13'b1000100000110,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110101,
13'b1000101110110,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1011101000101,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101110100,
13'b1100100100100,
13'b1100100110100,
13'b1100100110101,
13'b1100101000100,
13'b1100101000101,
13'b1100101010100: edge_mask_reg_512p1[363] <= 1'b1;
 		default: edge_mask_reg_512p1[363] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001001001,
13'b100001011010,
13'b101000111000,
13'b101000111001,
13'b101001001001,
13'b101001001010,
13'b101001011010,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b111000111001,
13'b111000111010,
13'b1010000010111,
13'b1010000011000,
13'b1011000010110,
13'b1011000010111,
13'b1100000010110,
13'b1100000010111: edge_mask_reg_512p1[364] <= 1'b1;
 		default: edge_mask_reg_512p1[364] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001001001,
13'b101000111000,
13'b101000111001,
13'b101001001001,
13'b101001001010,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b111000111001,
13'b111000111010,
13'b1010000010111,
13'b1010000011000,
13'b1011000010110,
13'b1011000010111,
13'b1100000010110,
13'b1100000010111: edge_mask_reg_512p1[365] <= 1'b1;
 		default: edge_mask_reg_512p1[365] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101010,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b111100001010,
13'b111100001011,
13'b111100011010,
13'b111100011011,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111000,
13'b111101111010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1000101101001,
13'b1000101111000,
13'b1001100100111,
13'b1001100101000,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101111000,
13'b1010100100111,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101111000,
13'b1011100100111,
13'b1011100101000,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1011101101000,
13'b1011101110111,
13'b1100100100111,
13'b1100100101000,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110111,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1110101100110,
13'b1110101100111,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111,
13'b1111101100110,
13'b1111101100111: edge_mask_reg_512p1[366] <= 1'b1;
 		default: edge_mask_reg_512p1[366] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101010,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b111100001010,
13'b111100001011,
13'b111100011010,
13'b111100011011,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111000,
13'b111101111010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1000101101001,
13'b1000101111000,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101111000,
13'b1010100100111,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101111000,
13'b1011100100111,
13'b1011100101000,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1011101101000,
13'b1011101110111,
13'b1100100100111,
13'b1100100101000,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110111,
13'b1101100100111,
13'b1101100101000,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1110101100110,
13'b1110101100111,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111,
13'b1111101100110,
13'b1111101100111: edge_mask_reg_512p1[367] <= 1'b1;
 		default: edge_mask_reg_512p1[367] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001001001,
13'b101000111001,
13'b101001001001,
13'b101001001010,
13'b110000111001,
13'b110000111010,
13'b110001001010,
13'b1010000010111,
13'b1011000010110,
13'b1011000010111,
13'b1100000010110,
13'b1100000010111: edge_mask_reg_512p1[368] <= 1'b1;
 		default: edge_mask_reg_512p1[368] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001111001,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111010,
13'b11001111011,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111010,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000111,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001011001,
13'b111001011010,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000001000110,
13'b1000001000111,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000110,
13'b1001001000111,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000110,
13'b1010001000111,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1100000010101,
13'b1100000010110,
13'b1100000010111,
13'b1100000100101,
13'b1100000100110,
13'b1100000110101,
13'b1101000010101,
13'b1101000010110,
13'b1101000100101,
13'b1101000100110: edge_mask_reg_512p1[369] <= 1'b1;
 		default: edge_mask_reg_512p1[369] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10001101000,
13'b10001101001,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101001,
13'b101001101010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011001,
13'b110001011010,
13'b110001101010,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001001001,
13'b111001001010,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000110110,
13'b1000000110111,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1010000010111,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1011000010110,
13'b1011000010111,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110110,
13'b1100000010101,
13'b1100000010110,
13'b1100000010111,
13'b1100000100100,
13'b1100000100101,
13'b1100000100110,
13'b1100000100111,
13'b1101000010101,
13'b1101000010110,
13'b1101000100101: edge_mask_reg_512p1[370] <= 1'b1;
 		default: edge_mask_reg_512p1[370] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011010,
13'b11110011011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b100110011011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110011011,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011010,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111010,
13'b111101111011,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1001100000111,
13'b1001100001000,
13'b1001100010111,
13'b1001100011000,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1010100000111,
13'b1010100001000,
13'b1010100010111,
13'b1010100011000,
13'b1010100100111,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1011100000111,
13'b1011100001000,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1011101101000,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1100101101000,
13'b1101100010110,
13'b1101100010111,
13'b1101100011000,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1110100010110,
13'b1110100100110,
13'b1110100100111,
13'b1110100110110,
13'b1110100110111,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1110101100110,
13'b1111100100110,
13'b1111100110110,
13'b1111100110111,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111: edge_mask_reg_512p1[371] <= 1'b1;
 		default: edge_mask_reg_512p1[371] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b100110011011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110011011,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011010,
13'b110110011011,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1001100000111,
13'b1001100001000,
13'b1001100010111,
13'b1001100011000,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1010100000111,
13'b1010100001000,
13'b1010100010111,
13'b1010100011000,
13'b1010100100111,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1011100000111,
13'b1011100001000,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1011101101000,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1100101101000,
13'b1101100010110,
13'b1101100010111,
13'b1101100011000,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1110100010110,
13'b1110100100110,
13'b1110100100111,
13'b1110100110110,
13'b1110100110111,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1110101100110,
13'b1111100100110,
13'b1111100110110,
13'b1111100110111,
13'b1111101000110,
13'b1111101000111,
13'b1111101010111: edge_mask_reg_512p1[372] <= 1'b1;
 		default: edge_mask_reg_512p1[372] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111011,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101010,
13'b11101101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101010,
13'b100101101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101010,
13'b101101101011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111001,
13'b111100111010,
13'b111101001010,
13'b111101001011,
13'b1000011100111,
13'b1000011101000,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1001011100111,
13'b1001011101000,
13'b1001011110111,
13'b1001011111000,
13'b1001011111001,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100010111,
13'b1001100011000,
13'b1001100011001,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1010011010111,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010011111001,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100001001,
13'b1010100010111,
13'b1010100011000,
13'b1010100011001,
13'b1010100100111,
13'b1010100101000,
13'b1011011100110,
13'b1011011100111,
13'b1011011101000,
13'b1011011110110,
13'b1011011110111,
13'b1011011111000,
13'b1011100000110,
13'b1011100000111,
13'b1011100001000,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100100111,
13'b1011100101000,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100011111000,
13'b1100100000110,
13'b1100100000111,
13'b1100100001000,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1100100100111,
13'b1100100101000,
13'b1101011100110,
13'b1101011100111,
13'b1101011110110,
13'b1101011110111,
13'b1101011111000,
13'b1101100000110,
13'b1101100000111,
13'b1101100001000,
13'b1101100010110,
13'b1101100010111,
13'b1101100011000,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1110011110110,
13'b1110011110111,
13'b1110100000110,
13'b1110100000111,
13'b1110100010110,
13'b1110100010111,
13'b1111100000110,
13'b1111100000111,
13'b1111100010110,
13'b1111100010111: edge_mask_reg_512p1[373] <= 1'b1;
 		default: edge_mask_reg_512p1[373] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b101111001001,
13'b101111001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b111110101010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100,
13'b1011110000100,
13'b1011110010100: edge_mask_reg_512p1[374] <= 1'b1;
 		default: edge_mask_reg_512p1[374] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100001001,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b101111001001,
13'b101111001010,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b111110101010,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1010101000100,
13'b1010101000101,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100,
13'b1011110000100,
13'b1011110010100: edge_mask_reg_512p1[375] <= 1'b1;
 		default: edge_mask_reg_512p1[375] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b101111001001,
13'b101111001010,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b111110101010,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1010101000100,
13'b1010101000101,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011110000100,
13'b1011110010100,
13'b1100101010100,
13'b1100101100100: edge_mask_reg_512p1[376] <= 1'b1;
 		default: edge_mask_reg_512p1[376] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111010,
13'b11101111011,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b110011001001,
13'b110011001010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1001011100101,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000101,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010101000101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011101000101,
13'b1100100000100,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100110101,
13'b1100101000101: edge_mask_reg_512p1[377] <= 1'b1;
 		default: edge_mask_reg_512p1[377] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111010,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111010,
13'b110001101010,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b111001111010,
13'b111001111011,
13'b111010001010,
13'b111010001011,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b1000010011000,
13'b1000010011001,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011011010,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1001010011000,
13'b1001010011001,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011100111,
13'b1001011101000,
13'b1001011101001,
13'b1001011110111,
13'b1001011111000,
13'b1010010010111,
13'b1010010011000,
13'b1010010100111,
13'b1010010101000,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110111,
13'b1010011111000,
13'b1011010010111,
13'b1011010011000,
13'b1011010100111,
13'b1011010101000,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100110,
13'b1011011100111,
13'b1011011101000,
13'b1011011110110,
13'b1011011110111,
13'b1011011111000,
13'b1100010010111,
13'b1100010011000,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1100011110110,
13'b1100011110111,
13'b1100011111000,
13'b1101010010111,
13'b1101010011000,
13'b1101010100111,
13'b1101010101000,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1101011100110,
13'b1101011100111,
13'b1101011101000,
13'b1101011110110,
13'b1101011110111,
13'b1110010110110,
13'b1110010110111,
13'b1110011000110,
13'b1110011000111,
13'b1110011010110,
13'b1110011010111,
13'b1110011100110,
13'b1110011100111,
13'b1110011110110,
13'b1111010110110,
13'b1111010110111,
13'b1111011000110,
13'b1111011000111,
13'b1111011010110: edge_mask_reg_512p1[378] <= 1'b1;
 		default: edge_mask_reg_512p1[378] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111110111011,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111001011,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111011011,
13'b111111100111,
13'b111111101000,
13'b1000110010111,
13'b1000110011000,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000110111010,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111001010,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111100110,
13'b1001111100111,
13'b1010110010110,
13'b1010110010111,
13'b1010110100110,
13'b1010110100111,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100110,
13'b1010111100111,
13'b1011110010110,
13'b1011110010111,
13'b1011110100110,
13'b1011110100111,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100110,
13'b1011111100111,
13'b1100110100110,
13'b1100110100111,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111010101,
13'b1100111010110,
13'b1101110100110,
13'b1101110110101,
13'b1101110110110,
13'b1101111000101,
13'b1101111000110,
13'b1101111010101,
13'b1101111010110,
13'b1110110100110,
13'b1110110110110,
13'b1110111000110: edge_mask_reg_512p1[379] <= 1'b1;
 		default: edge_mask_reg_512p1[379] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111110111011,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111001011,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111011011,
13'b111111100111,
13'b111111101000,
13'b1000110010111,
13'b1000110011000,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000110111010,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111001010,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111100110,
13'b1001111100111,
13'b1010110010110,
13'b1010110010111,
13'b1010110100110,
13'b1010110100111,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1011110010110,
13'b1011110010111,
13'b1011110100110,
13'b1011110100111,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1100110100110,
13'b1100110100111,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111010101,
13'b1100111010110,
13'b1100111100101,
13'b1100111100110,
13'b1101110100110,
13'b1101110110101,
13'b1101110110110,
13'b1101111000101,
13'b1101111000110,
13'b1101111010101,
13'b1101111010110,
13'b1101111100101,
13'b1110110100110,
13'b1110110110110,
13'b1110111000110: edge_mask_reg_512p1[380] <= 1'b1;
 		default: edge_mask_reg_512p1[380] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111110111011,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111001011,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111011011,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000110010111,
13'b1000110011000,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000110111010,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111001010,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111011010,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010110010110,
13'b1010110010111,
13'b1010110100110,
13'b1010110100111,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1011110010110,
13'b1011110010111,
13'b1011110100110,
13'b1011110100111,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110110,
13'b1011111110111,
13'b1100110100110,
13'b1100110100111,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111010101,
13'b1100111010110,
13'b1100111010111,
13'b1100111100101,
13'b1100111100110,
13'b1101110100110,
13'b1101110110101,
13'b1101110110110,
13'b1101111000101,
13'b1101111000110,
13'b1101111010101,
13'b1101111010110,
13'b1101111100101,
13'b1101111100110,
13'b1110110100110,
13'b1110110110110,
13'b1110111000110: edge_mask_reg_512p1[381] <= 1'b1;
 		default: edge_mask_reg_512p1[381] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011010,
13'b11010011011,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011010,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100111,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001111001,
13'b111001111010,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001100110,
13'b1000001100111,
13'b1001000100110,
13'b1001000100111,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010110,
13'b1001001010111,
13'b1001001100110,
13'b1001001100111,
13'b1010000010111,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001010110,
13'b1010001010111,
13'b1010001100110,
13'b1010001100111,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1011001000101,
13'b1011001000110,
13'b1011001000111,
13'b1011001010110,
13'b1011001010111,
13'b1011001100110,
13'b1011001100111,
13'b1100000010101,
13'b1100000010110,
13'b1100000100101,
13'b1100000100110,
13'b1100000110101,
13'b1100000110110,
13'b1100001000101,
13'b1100001000110,
13'b1101000010101,
13'b1101000010110,
13'b1101000100101,
13'b1101000100110,
13'b1101000110101,
13'b1101000110110,
13'b1101001000101: edge_mask_reg_512p1[382] <= 1'b1;
 		default: edge_mask_reg_512p1[382] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111010,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111001,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b110011011001,
13'b110011011010,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101010011,
13'b1000101010100,
13'b1001011110101,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010100,
13'b1011100000100,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100: edge_mask_reg_512p1[383] <= 1'b1;
 		default: edge_mask_reg_512p1[383] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101110101000,
13'b101110101001,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110111000,
13'b111111000110,
13'b111111001000,
13'b111111001001,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000111000101,
13'b1000111000110,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100110,
13'b1000111100111,
13'b1001111000101,
13'b1001111000110,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010111000101,
13'b1010111000110,
13'b1010111010101,
13'b1010111010110,
13'b1010111100101,
13'b1010111100110,
13'b1011111000101,
13'b1011111000110,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1100111000101,
13'b1100111010100,
13'b1100111010101,
13'b1100111010110,
13'b1100111100100,
13'b1100111100101,
13'b1100111100110,
13'b1100111110101,
13'b1100111110110,
13'b1101111010100,
13'b1101111010101,
13'b1101111100100,
13'b1101111100101,
13'b1101111110101,
13'b1110111010100,
13'b1110111100100: edge_mask_reg_512p1[384] <= 1'b1;
 		default: edge_mask_reg_512p1[384] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000100,
13'b11101000101,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b101010011001,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110010101001,
13'b110010101010,
13'b110010110100,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b1000011010011,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1001011100011,
13'b1001011110011,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100110011: edge_mask_reg_512p1[385] <= 1'b1;
 		default: edge_mask_reg_512p1[385] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001010,
13'b11110001011,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101010100,
13'b1001101010101,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010100,
13'b1010101010101,
13'b1011100010110,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010100,
13'b1011101010101,
13'b1100100100110,
13'b1100100100111,
13'b1100100110100,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010101,
13'b1101101010110: edge_mask_reg_512p1[386] <= 1'b1;
 		default: edge_mask_reg_512p1[386] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100101010,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010101,
13'b10101010110,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001010,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101011001,
13'b111101011010,
13'b111101100011,
13'b111101101001,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101100011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100: edge_mask_reg_512p1[387] <= 1'b1;
 		default: edge_mask_reg_512p1[387] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1101001010,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011001,
13'b100110011010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110101,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110101,
13'b1010100100011,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101110100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[388] <= 1'b1;
 		default: edge_mask_reg_512p1[388] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1101001010,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b101110011010,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110101,
13'b1000101110110,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110101,
13'b1010100100011,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[389] <= 1'b1;
 		default: edge_mask_reg_512p1[389] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111010,
13'b11101111011,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111010,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b111011011010,
13'b111011011011,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b1000011111000,
13'b1000011111001,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100011010,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100101010,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101001000,
13'b1001011111000,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100010111,
13'b1001100011000,
13'b1001100011001,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101001000,
13'b1010011110111,
13'b1010011111000,
13'b1010100000111,
13'b1010100001000,
13'b1010100010111,
13'b1010100011000,
13'b1010100100111,
13'b1010100101000,
13'b1010100101001,
13'b1010100110111,
13'b1010100111000,
13'b1010101001000,
13'b1011011110111,
13'b1011011111000,
13'b1011100000111,
13'b1011100001000,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1100011110111,
13'b1100011111000,
13'b1100100000111,
13'b1100100001000,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1101100000111,
13'b1101100001000,
13'b1101100010110,
13'b1101100010111,
13'b1101100011000,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1110100010110,
13'b1110100010111,
13'b1110100100110,
13'b1110100100111,
13'b1110100110110,
13'b1111100100110: edge_mask_reg_512p1[390] <= 1'b1;
 		default: edge_mask_reg_512p1[390] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100: edge_mask_reg_512p1[391] <= 1'b1;
 		default: edge_mask_reg_512p1[391] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100: edge_mask_reg_512p1[392] <= 1'b1;
 		default: edge_mask_reg_512p1[392] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101001,
13'b11101101010,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010011,
13'b101101010100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000011,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101001001,
13'b1000011000101,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001101000011,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100: edge_mask_reg_512p1[393] <= 1'b1;
 		default: edge_mask_reg_512p1[393] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101001,
13'b11101101010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010011,
13'b101101010100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110010101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000011,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101001001,
13'b1000011000101,
13'b1000011010100,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1001011010100,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1011011110100,
13'b1011100000100: edge_mask_reg_512p1[394] <= 1'b1;
 		default: edge_mask_reg_512p1[394] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011001,
13'b101011011010,
13'b110000110110,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b111000110101,
13'b111000110110,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b1000000110101,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100101,
13'b1000010100110,
13'b1000010110101,
13'b1001001000101,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100101,
13'b1001010100110,
13'b1010001010100,
13'b1010001010101,
13'b1010001100100,
13'b1010001100101,
13'b1010001110100,
13'b1010001110101,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1011001010100,
13'b1011001100100,
13'b1011001110100,
13'b1011010000100,
13'b1011010010100: edge_mask_reg_512p1[395] <= 1'b1;
 		default: edge_mask_reg_512p1[395] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011010,
13'b10011011011,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001001,
13'b101011001010,
13'b110000110110,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b111000110101,
13'b111000110110,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b1000000110101,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100101,
13'b1000010100110,
13'b1001001000101,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100101,
13'b1001010100110,
13'b1010001010100,
13'b1010001010101,
13'b1010001100100,
13'b1010001100101,
13'b1010001110100,
13'b1010001110101,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1011001010100,
13'b1011001100100,
13'b1011001100101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101: edge_mask_reg_512p1[396] <= 1'b1;
 		default: edge_mask_reg_512p1[396] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b110001101001,
13'b110001101010,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1001010000101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1011010010100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[397] <= 1'b1;
 		default: edge_mask_reg_512p1[397] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010111001,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b101001011001,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b110001101001,
13'b110001101010,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100100,
13'b1000011100101,
13'b1001010000100,
13'b1001010000101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1010010000100,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1011010010100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[398] <= 1'b1;
 		default: edge_mask_reg_512p1[398] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010111,
13'b1000101011000,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1011100010110,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100101,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010101,
13'b1101101010110,
13'b1101101100101,
13'b1110100110101,
13'b1110100110110,
13'b1110101000101,
13'b1110101000110,
13'b1110101010101,
13'b1110101010110: edge_mask_reg_512p1[399] <= 1'b1;
 		default: edge_mask_reg_512p1[399] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010111,
13'b1000101011000,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010110,
13'b1010101010111,
13'b1011100010110,
13'b1011100010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100101,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010101,
13'b1101101010110,
13'b1101101100101,
13'b1110100110101,
13'b1110100110110,
13'b1110101000101,
13'b1110101000110,
13'b1110101010101,
13'b1110101010110: edge_mask_reg_512p1[400] <= 1'b1;
 		default: edge_mask_reg_512p1[400] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100010110,
13'b1000100010111,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111010,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010111,
13'b1000101011000,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010110,
13'b1010101010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100101,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010101,
13'b1101101010110,
13'b1101101100101,
13'b1110100110110,
13'b1110101000101,
13'b1110101000110,
13'b1110101010101,
13'b1110101010110: edge_mask_reg_512p1[401] <= 1'b1;
 		default: edge_mask_reg_512p1[401] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010110,
13'b110101010111,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100000101,
13'b1000100000110,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010101,
13'b1000101010110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010101,
13'b1001101010110,
13'b1010100010100,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101010101,
13'b1010101010110,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1011101000101,
13'b1011101010100,
13'b1011101010101,
13'b1100100100100,
13'b1100100110100,
13'b1100100110101,
13'b1100101000100,
13'b1100101000101: edge_mask_reg_512p1[402] <= 1'b1;
 		default: edge_mask_reg_512p1[402] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b110110001010,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100101,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010100,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100: edge_mask_reg_512p1[403] <= 1'b1;
 		default: edge_mask_reg_512p1[403] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010110,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b111110101010,
13'b1000100110101,
13'b1000100110110,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1001110000110,
13'b1001110010101,
13'b1001110010110,
13'b1010101000100,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010101,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1100101010100,
13'b1100101100100,
13'b1100101100101,
13'b1100101110100,
13'b1100101110101,
13'b1100110000100,
13'b1100110000101: edge_mask_reg_512p1[404] <= 1'b1;
 		default: edge_mask_reg_512p1[404] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010110,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b111110101010,
13'b1000100110101,
13'b1000100110110,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1001100110101,
13'b1001100110110,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010101,
13'b1001110010110,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010101,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1100101010100,
13'b1100101100100,
13'b1100101100101,
13'b1100101110100,
13'b1100101110101,
13'b1100110000100,
13'b1100110000101: edge_mask_reg_512p1[405] <= 1'b1;
 		default: edge_mask_reg_512p1[405] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110101001,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010011,
13'b1001110010100,
13'b1001110100011,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010110000011,
13'b1010110000100,
13'b1010110010011,
13'b1010110010100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[406] <= 1'b1;
 		default: edge_mask_reg_512p1[406] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100001001,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110101001,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010011,
13'b1001110010100,
13'b1001110100011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000011,
13'b1010110000100,
13'b1010110010011,
13'b1010110010100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[407] <= 1'b1;
 		default: edge_mask_reg_512p1[407] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101001,
13'b11110101010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1001100110100,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100,
13'b1100101000100,
13'b1100101010100: edge_mask_reg_512p1[408] <= 1'b1;
 		default: edge_mask_reg_512p1[408] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000110,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000101,
13'b1000110000110,
13'b1001100110100,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101110100,
13'b1100101000100,
13'b1100101010100,
13'b1100101100100: edge_mask_reg_512p1[409] <= 1'b1;
 		default: edge_mask_reg_512p1[409] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b111110011010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1001100110100,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1100101000100,
13'b1100101010100,
13'b1100101100100: edge_mask_reg_512p1[410] <= 1'b1;
 		default: edge_mask_reg_512p1[410] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b110010011001,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011101100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110011111100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100001100,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100011100,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011010,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1010011000101,
13'b1010011000110,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1011011010101,
13'b1011011010110,
13'b1011011100101,
13'b1011011100110,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010101,
13'b1011100010110,
13'b1011100100101,
13'b1011100100110,
13'b1100011010101,
13'b1100011100101,
13'b1100011100110,
13'b1100011110101,
13'b1100011110110,
13'b1100100000101,
13'b1100100000110,
13'b1100100010101,
13'b1100100010110,
13'b1100100100101,
13'b1100100100110,
13'b1101011100101,
13'b1101011110101,
13'b1101011110110,
13'b1101100000101,
13'b1101100000110,
13'b1101100010101,
13'b1101100010110,
13'b1101100100110: edge_mask_reg_512p1[411] <= 1'b1;
 		default: edge_mask_reg_512p1[411] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100101010,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010111,
13'b1000101011000,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010110,
13'b1010101010111,
13'b1011100010110,
13'b1011100010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1100100010111,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100101,
13'b1101100100110,
13'b1101100100111,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101010101,
13'b1101101010110,
13'b1101101100101,
13'b1110100110110,
13'b1110100110111,
13'b1110101000101,
13'b1110101000110,
13'b1110101000111,
13'b1110101010101,
13'b1110101010110,
13'b1111100110110: edge_mask_reg_512p1[412] <= 1'b1;
 		default: edge_mask_reg_512p1[412] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110001001,
13'b111110011001,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000101,
13'b1000110000110,
13'b1001100110100,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1100101000100,
13'b1100101010100,
13'b1100101100100,
13'b1100101110100: edge_mask_reg_512p1[413] <= 1'b1;
 		default: edge_mask_reg_512p1[413] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001000,
13'b100111001001,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100110,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100101,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100101,
13'b1010101000100,
13'b1010101000101,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1011110010100,
13'b1100101010100,
13'b1100101100100,
13'b1100101110100,
13'b1100110000100: edge_mask_reg_512p1[414] <= 1'b1;
 		default: edge_mask_reg_512p1[414] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001000,
13'b100111001001,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100110,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100101,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100101,
13'b1010101000100,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1011110010100,
13'b1100101100100,
13'b1100101110100,
13'b1100110000100: edge_mask_reg_512p1[415] <= 1'b1;
 		default: edge_mask_reg_512p1[415] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011010,
13'b11110011011,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b101011001010,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101001,
13'b111101101010,
13'b111101111010,
13'b1000011110111,
13'b1000011111000,
13'b1000100000111,
13'b1000100001000,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1001011110111,
13'b1001011111000,
13'b1001100000111,
13'b1001100001000,
13'b1001100010111,
13'b1001100011000,
13'b1001100100111,
13'b1001100101000,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101101000,
13'b1010011110111,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101010111,
13'b1010101011000,
13'b1011011110111,
13'b1011100000110,
13'b1011100000111,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1100011110111,
13'b1100100000110,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1101100000111,
13'b1101100010110,
13'b1101100010111,
13'b1101100100110,
13'b1101100100111,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1110100010110,
13'b1110100100110,
13'b1110100100111,
13'b1110100110110,
13'b1110100110111,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1111100100110,
13'b1111100110110,
13'b1111101000110,
13'b1111101010110: edge_mask_reg_512p1[416] <= 1'b1;
 		default: edge_mask_reg_512p1[416] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011010,
13'b11110011011,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b100110011011,
13'b101011001010,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110011011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111010,
13'b111101111011,
13'b1000011110111,
13'b1000011111000,
13'b1000100000111,
13'b1000100001000,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1001011110111,
13'b1001011111000,
13'b1001100000111,
13'b1001100001000,
13'b1001100010111,
13'b1001100011000,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1010011110111,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101101000,
13'b1011011110111,
13'b1011100000110,
13'b1011100000111,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1100011110111,
13'b1100100000110,
13'b1100100000111,
13'b1100100010110,
13'b1100100010111,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1101100000111,
13'b1101100010110,
13'b1101100010111,
13'b1101100100110,
13'b1101100100111,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1110100010110,
13'b1110100100110,
13'b1110100100111,
13'b1110100110110,
13'b1110100110111,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1111100100110,
13'b1111100110110,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111: edge_mask_reg_512p1[417] <= 1'b1;
 		default: edge_mask_reg_512p1[417] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001011,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100001100,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100011100,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100101100,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110100111100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111010,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000101,
13'b1001101000110,
13'b1010100000110,
13'b1010100000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000101,
13'b1010101000110,
13'b1011100010110,
13'b1011100010111,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101010101,
13'b1100100010111,
13'b1100100100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100101000101,
13'b1100101000110,
13'b1101100100101,
13'b1101100100110,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110: edge_mask_reg_512p1[418] <= 1'b1;
 		default: edge_mask_reg_512p1[418] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001010,
13'b10110001011,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100001100,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100011100,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100101100,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110100111100,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b111101101010,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000101,
13'b1001101000110,
13'b1010100000110,
13'b1010100000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000101,
13'b1010101000110,
13'b1011100010110,
13'b1011100010111,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101010101,
13'b1100100010111,
13'b1100100100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100101000101,
13'b1100101000110,
13'b1100101010101,
13'b1101100100101,
13'b1101100100110,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110: edge_mask_reg_512p1[419] <= 1'b1;
 		default: edge_mask_reg_512p1[419] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110100,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110011,
13'b101101110100,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110011,
13'b110101110100,
13'b110101111000,
13'b110101111001,
13'b111011100100,
13'b111011101001,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101011000,
13'b111101011001,
13'b111101100011,
13'b111101101000,
13'b111101101001,
13'b1000011110011,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101000100,
13'b1000101010011,
13'b1000101100011,
13'b1001100000011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001101000011,
13'b1010100010011,
13'b1010100100011,
13'b1010100110011: edge_mask_reg_512p1[420] <= 1'b1;
 		default: edge_mask_reg_512p1[420] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001010,
13'b10010001011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001010,
13'b11010001011,
13'b100001001000,
13'b100001001001,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001010,
13'b100010001011,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001010,
13'b101010001011,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111010,
13'b110001111011,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111000111011,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001001011,
13'b111001011010,
13'b111001011011,
13'b111001101010,
13'b111001101011,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000101010,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000000111010,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110110,
13'b1001000110111,
13'b1001000111000,
13'b1001001000110,
13'b1001001000111,
13'b1001001001000,
13'b1010000010111,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000110,
13'b1010001000111,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1011001000110,
13'b1011001000111,
13'b1100000010101,
13'b1100000010110,
13'b1100000010111,
13'b1100000100101,
13'b1100000100110,
13'b1100000100111,
13'b1100000110101,
13'b1100000110110,
13'b1101000010101,
13'b1101000010110,
13'b1101000100101,
13'b1101000100110,
13'b1101000110110: edge_mask_reg_512p1[421] <= 1'b1;
 		default: edge_mask_reg_512p1[421] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000101,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111001,
13'b100101111010,
13'b101011011001,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101010011,
13'b111101010100,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100: edge_mask_reg_512p1[422] <= 1'b1;
 		default: edge_mask_reg_512p1[422] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000101,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001010,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001001,
13'b100110001010,
13'b101011011001,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100: edge_mask_reg_512p1[423] <= 1'b1;
 		default: edge_mask_reg_512p1[423] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010101,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010011,
13'b100101010100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b101011011001,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010011,
13'b101101010100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b111011111001,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101010010,
13'b111101010011,
13'b111101011001,
13'b111101100011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101010011,
13'b1000101100011,
13'b1001100010011,
13'b1001100100011,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011: edge_mask_reg_512p1[424] <= 1'b1;
 		default: edge_mask_reg_512p1[424] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011010,
13'b11100011011,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001001010,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011010,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010001100,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010011100,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010101100,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011001100,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b111001101010,
13'b111001101011,
13'b111001111010,
13'b111001111011,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101000,
13'b111011101010,
13'b111011101011,
13'b111011111010,
13'b111011111011,
13'b1000001111000,
13'b1000010000111,
13'b1000010001000,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010011010,
13'b1000010011011,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010101010,
13'b1000010101011,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011101000,
13'b1001010000111,
13'b1001010001000,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010111,
13'b1001011011000,
13'b1001011101000,
13'b1010010000110,
13'b1010010000111,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1011010000111,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100110,
13'b1100010010110,
13'b1100010010111,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100110,
13'b1101010100110,
13'b1101010110110,
13'b1101010110111,
13'b1101011000110,
13'b1101011000111,
13'b1101011010110,
13'b1101011010111,
13'b1101011100110,
13'b1110010110110,
13'b1110011000110,
13'b1110011010110: edge_mask_reg_512p1[425] <= 1'b1;
 		default: edge_mask_reg_512p1[425] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000011110101,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1001011110101,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000101,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010101000100,
13'b1010101000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1011101000101,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100110100,
13'b1100100110101: edge_mask_reg_512p1[426] <= 1'b1;
 		default: edge_mask_reg_512p1[426] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111010,
13'b11101111011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b1000011110101,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1001011110101,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000101,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010101000100,
13'b1010101000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011101000100,
13'b1011101000101,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100110100,
13'b1100100110101,
13'b1100101000101: edge_mask_reg_512p1[427] <= 1'b1;
 		default: edge_mask_reg_512p1[427] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111010,
13'b11100111011,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b110010011001,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000101,
13'b1010011000101,
13'b1010011000110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011011010101,
13'b1011011010110,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000101,
13'b1101011100101: edge_mask_reg_512p1[428] <= 1'b1;
 		default: edge_mask_reg_512p1[428] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111010,
13'b11100111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b101010001010,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000101,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011011000110,
13'b1011011010101,
13'b1011011010110,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1100011010101,
13'b1100011010110,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000101,
13'b1101011100101,
13'b1101011110101: edge_mask_reg_512p1[429] <= 1'b1;
 		default: edge_mask_reg_512p1[429] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1010100110101,
13'b1011011110101,
13'b1011011110110,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1100100000100,
13'b1100100000101,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1101100010101: edge_mask_reg_512p1[430] <= 1'b1;
 		default: edge_mask_reg_512p1[430] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101010,
13'b111100001010,
13'b111100001011,
13'b111100011010,
13'b111100011011,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b1000100101000,
13'b1000100101001,
13'b1000100111000,
13'b1000100111001,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1000101101001,
13'b1000101111000,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1001101101001,
13'b1001101111000,
13'b1010100100111,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101111000,
13'b1011100100111,
13'b1011100101000,
13'b1011100110111,
13'b1011100111000,
13'b1011101000111,
13'b1011101001000,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1011101111000,
13'b1100100100111,
13'b1100100101000,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1100101101000,
13'b1100101110111,
13'b1100101111000,
13'b1101100100111,
13'b1101100101000,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110111,
13'b1101101111000,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1111101000111,
13'b1111101010111,
13'b1111101100111: edge_mask_reg_512p1[431] <= 1'b1;
 		default: edge_mask_reg_512p1[431] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101010,
13'b111100001010,
13'b111100011010,
13'b111100011011,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b1000100111000,
13'b1000100111001,
13'b1000101001000,
13'b1000101001001,
13'b1000101011000,
13'b1000101011001,
13'b1000101101000,
13'b1000101101001,
13'b1000101111000,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101011000,
13'b1001101011001,
13'b1001101101000,
13'b1001101101001,
13'b1001101111000,
13'b1010100101000,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101111000,
13'b1011100101000,
13'b1011100110111,
13'b1011100111000,
13'b1011101000111,
13'b1011101001000,
13'b1011101010111,
13'b1011101011000,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1011101111000,
13'b1100100101000,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100111,
13'b1100101101000,
13'b1100101110111,
13'b1100101111000,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110111,
13'b1101101111000,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1111101000111,
13'b1111101010111,
13'b1111101100111: edge_mask_reg_512p1[432] <= 1'b1;
 		default: edge_mask_reg_512p1[432] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001001,
13'b100100001010,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011101001,
13'b111011101010,
13'b1000001110101,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1001010000101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010101,
13'b1010010010011,
13'b1010010010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1011010010100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[433] <= 1'b1;
 		default: edge_mask_reg_512p1[433] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001010,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011101001,
13'b1000001110101,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1001010000101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000100,
13'b1001011000101,
13'b1001011010101,
13'b1010010010011,
13'b1010010010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000100,
13'b1011010010100,
13'b1011010100100,
13'b1011010110100,
13'b1011011000100: edge_mask_reg_512p1[434] <= 1'b1;
 		default: edge_mask_reg_512p1[434] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011001,
13'b11100011010,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011001,
13'b100100011010,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001001,
13'b110100001010,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001001,
13'b111010001010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b1000001110101,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1001010010011,
13'b1001010010100,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100101,
13'b1010010010100,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100: edge_mask_reg_512p1[435] <= 1'b1;
 		default: edge_mask_reg_512p1[435] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101001001,
13'b111101001010,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110100,
13'b1000100110101,
13'b1001011110101,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001101000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000100,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100110100,
13'b1100100110101: edge_mask_reg_512p1[436] <= 1'b1;
 		default: edge_mask_reg_512p1[436] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101010,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110100,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b101011101000,
13'b101011101001,
13'b101011110100,
13'b101011110101,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110011,
13'b101101110100,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b110011110100,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101101000,
13'b110101101001,
13'b110101110011,
13'b110101110100,
13'b110101111000,
13'b110101111001,
13'b111011110100,
13'b111011111000,
13'b111011111001,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101011000,
13'b111101011001,
13'b111101100011,
13'b111101101000,
13'b111101101001,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101000100,
13'b1000101010011,
13'b1000101100011,
13'b1001100010011,
13'b1001100100011,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101010011,
13'b1010100100011,
13'b1010100110011,
13'b1010101000011,
13'b1010101010011: edge_mask_reg_512p1[437] <= 1'b1;
 		default: edge_mask_reg_512p1[437] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101010,
13'b111011000100,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1001100110101,
13'b1010011110100,
13'b1010100000100,
13'b1010100010100,
13'b1010100010101,
13'b1010100100100,
13'b1010100110100,
13'b1011100010100: edge_mask_reg_512p1[438] <= 1'b1;
 		default: edge_mask_reg_512p1[438] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b101010101001,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101010,
13'b111011000100,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b1000011010011,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1001100110101,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1010100100100,
13'b1010100110100,
13'b1011100010100: edge_mask_reg_512p1[439] <= 1'b1;
 		default: edge_mask_reg_512p1[439] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101011010,
13'b1000011100101,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100110100,
13'b1011100110101,
13'b1100100010101,
13'b1100100100101,
13'b1100100110101: edge_mask_reg_512p1[440] <= 1'b1;
 		default: edge_mask_reg_512p1[440] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101001010,
13'b111101011010,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100110100,
13'b1011100110101,
13'b1100100010101,
13'b1100100100101,
13'b1100100110101: edge_mask_reg_512p1[441] <= 1'b1;
 		default: edge_mask_reg_512p1[441] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101010,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100101100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110100111100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101001100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101011100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110110,
13'b110101110111,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011001,
13'b110110011010,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100111010,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001010,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110101,
13'b1000101110110,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110101,
13'b1001101110110,
13'b1010100110100,
13'b1010100110101,
13'b1010101000100,
13'b1010101000101,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1011101000101,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101: edge_mask_reg_512p1[442] <= 1'b1;
 		default: edge_mask_reg_512p1[442] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110111001,
13'b11110111010,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110011100,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110011100,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110101100,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010111,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111110111011,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111001011,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111011011,
13'b1000110010111,
13'b1000110011000,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000110111010,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111001001,
13'b1000111001010,
13'b1000111010111,
13'b1000111011000,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1010110010110,
13'b1010110010111,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110110,
13'b1010110110111,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111010110,
13'b1010111010111,
13'b1010111011000,
13'b1011110010110,
13'b1011110010111,
13'b1011110100110,
13'b1011110100111,
13'b1011110110110,
13'b1011110110111,
13'b1011111000110,
13'b1011111000111,
13'b1011111010110,
13'b1011111010111,
13'b1100110100110,
13'b1100110100111,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111010111,
13'b1101110100110,
13'b1101110110110,
13'b1101110110111,
13'b1101111000110,
13'b1101111000111,
13'b1110110100110,
13'b1110110110110,
13'b1110111000110,
13'b1111110110110,
13'b1111111000110: edge_mask_reg_512p1[443] <= 1'b1;
 		default: edge_mask_reg_512p1[443] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010100,
13'b1010100100100: edge_mask_reg_512p1[444] <= 1'b1;
 		default: edge_mask_reg_512p1[444] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010100,
13'b1010100100100: edge_mask_reg_512p1[445] <= 1'b1;
 		default: edge_mask_reg_512p1[445] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010100,
13'b1010100100100: edge_mask_reg_512p1[446] <= 1'b1;
 		default: edge_mask_reg_512p1[446] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000101,
13'b11011000110,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111011000100,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010100,
13'b1010100100100: edge_mask_reg_512p1[447] <= 1'b1;
 		default: edge_mask_reg_512p1[447] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000110,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110100,
13'b1001100110101,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1010100100100,
13'b1010100110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[448] <= 1'b1;
 		default: edge_mask_reg_512p1[448] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111001,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b100110011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101101100,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101101111100,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110011011,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100101100,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110100111100,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101001100,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101011100,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101101100,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011010,
13'b110110011011,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111010,
13'b111101111011,
13'b111110001010,
13'b111110001011,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111010,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101011010,
13'b1000101101000,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101100111,
13'b1001101101000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100110,
13'b1010101100111,
13'b1011100010110,
13'b1011100010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100101,
13'b1100101100110,
13'b1100101110110,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010110,
13'b1101101100110,
13'b1110100110110,
13'b1110101000110: edge_mask_reg_512p1[449] <= 1'b1;
 		default: edge_mask_reg_512p1[449] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001001001,
13'b110001001010,
13'b110001011001,
13'b110001011010,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011101001,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000100,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1011011000100,
13'b1100001110100,
13'b1100001110101,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101,
13'b1100010100100,
13'b1100010100101: edge_mask_reg_512p1[450] <= 1'b1;
 		default: edge_mask_reg_512p1[450] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001001001,
13'b110001001010,
13'b110001011001,
13'b110001011010,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000100,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1011011000100,
13'b1100001110100,
13'b1100001110101,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101,
13'b1100010100100,
13'b1100010100101: edge_mask_reg_512p1[451] <= 1'b1;
 		default: edge_mask_reg_512p1[451] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001001001,
13'b110001001010,
13'b110001011001,
13'b110001011010,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000101,
13'b1001011000110,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1100001110100,
13'b1100001110101,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101,
13'b1100010100100,
13'b1100010100101: edge_mask_reg_512p1[452] <= 1'b1;
 		default: edge_mask_reg_512p1[452] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001001001,
13'b110001001010,
13'b110001011001,
13'b110001011010,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011011001,
13'b111011011010,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000101,
13'b1000011000110,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000101,
13'b1001011000110,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1100001110100,
13'b1100001110101,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101,
13'b1100010100100,
13'b1100010100101: edge_mask_reg_512p1[453] <= 1'b1;
 		default: edge_mask_reg_512p1[453] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b1001111001,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b10001101000,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101010,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b110001001001,
13'b110001001010,
13'b110001011001,
13'b110001011010,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001001,
13'b110011001010,
13'b110011011001,
13'b110011011010,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011001001,
13'b111011001010,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110101,
13'b1000010110110,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110101,
13'b1001010110110,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1100001110100,
13'b1100001110101,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101: edge_mask_reg_512p1[454] <= 1'b1;
 		default: edge_mask_reg_512p1[454] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111010,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b100001001000,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b110001001001,
13'b110001001010,
13'b110001010110,
13'b110001011001,
13'b110001011010,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110101,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100101,
13'b1001010100110,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1100001110100,
13'b1100001110101,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101: edge_mask_reg_512p1[455] <= 1'b1;
 		default: edge_mask_reg_512p1[455] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111010,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b110000111001,
13'b110000111010,
13'b110001001001,
13'b110001001010,
13'b110001010101,
13'b110001010110,
13'b110001011001,
13'b110001011010,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100101,
13'b1001010100110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1011001100100,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1100001110100,
13'b1100001110101,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101: edge_mask_reg_512p1[456] <= 1'b1;
 		default: edge_mask_reg_512p1[456] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b110000111001,
13'b110000111010,
13'b110001000110,
13'b110001000111,
13'b110001001001,
13'b110001001010,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111001,
13'b110010111010,
13'b110011001001,
13'b110011001010,
13'b111000111001,
13'b111000111010,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b1000001000101,
13'b1000001000110,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100101,
13'b1001010100110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1011001010100,
13'b1011001010101,
13'b1011001100100,
13'b1011001100101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1100001100100,
13'b1100001100101,
13'b1100001110100,
13'b1100001110101,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101: edge_mask_reg_512p1[457] <= 1'b1;
 		default: edge_mask_reg_512p1[457] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101010,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001001,
13'b101111001010,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111001,
13'b110110111010,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110011010,
13'b111110101001,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1001100110101,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1010101000100,
13'b1010101010100,
13'b1010101010101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010100,
13'b1010110010101,
13'b1011101000100,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110010100,
13'b1100101100100,
13'b1100101110100,
13'b1100110000100: edge_mask_reg_512p1[458] <= 1'b1;
 		default: edge_mask_reg_512p1[458] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101001,
13'b1101101010,
13'b1101111010,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001000,
13'b100111001001,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100110,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b111101000101,
13'b111101000110,
13'b111101001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110001010,
13'b111110010101,
13'b111110010110,
13'b111110011001,
13'b111110101001,
13'b1000101000101,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100101,
13'b1001101000101,
13'b1001101010101,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1011101100100,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1011110010100,
13'b1100101110100,
13'b1100110000100: edge_mask_reg_512p1[459] <= 1'b1;
 		default: edge_mask_reg_512p1[459] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100010110,
13'b1000100010111,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111010,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010111,
13'b1000101011000,
13'b1001100010110,
13'b1001100010111,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1010100010110,
13'b1010100010111,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010110,
13'b1010101010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100101,
13'b1100101100110,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101010101,
13'b1101101010110,
13'b1101101100101,
13'b1101101100110,
13'b1110100110110,
13'b1110101000101,
13'b1110101000110,
13'b1110101010101,
13'b1110101010110,
13'b1110101100110,
13'b1111101000110: edge_mask_reg_512p1[460] <= 1'b1;
 		default: edge_mask_reg_512p1[460] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111001,
13'b1101111010,
13'b1110001010,
13'b1110011000,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001000,
13'b100111001001,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b110100111001,
13'b110100111010,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110110,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111001000,
13'b110111001001,
13'b111101001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110101001,
13'b111110111000,
13'b111110111001,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110101,
13'b1001101010100,
13'b1001101010101,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110101,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1011101100100,
13'b1011101110100,
13'b1011101110101,
13'b1011110000100,
13'b1011110000101,
13'b1011110010100,
13'b1011110100100,
13'b1100101110100,
13'b1100110000100: edge_mask_reg_512p1[461] <= 1'b1;
 		default: edge_mask_reg_512p1[461] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100111010,
13'b1101000101,
13'b1101000110,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010101,
13'b1101010110,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100101,
13'b1101100110,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110100,
13'b10101110101,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000100,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011001,
13'b11110011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000100,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b101011101000,
13'b101011101001,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110011,
13'b101101110100,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000011,
13'b101110000100,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011001,
13'b110011110100,
13'b110011111000,
13'b110011111001,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110011,
13'b110101110100,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100001001,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100010,
13'b111101100011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101110010,
13'b111101110011,
13'b111101111001,
13'b1000100010011,
13'b1000100100011,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101010011,
13'b1000101100011,
13'b1000101110011,
13'b1001100100011,
13'b1001100110011,
13'b1001101000011,
13'b1010100110011: edge_mask_reg_512p1[462] <= 1'b1;
 		default: edge_mask_reg_512p1[462] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000101,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110100,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110100,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101100100,
13'b111101101001,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101100011,
13'b1000101100100,
13'b1001100000011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100: edge_mask_reg_512p1[463] <= 1'b1;
 		default: edge_mask_reg_512p1[463] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000101,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110100,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110100,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101100100,
13'b111101101001,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101100011,
13'b1000101100100,
13'b1001100000011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1010100010011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100: edge_mask_reg_512p1[464] <= 1'b1;
 		default: edge_mask_reg_512p1[464] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000101,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110100,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110100,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101101001,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101100011,
13'b1000101100100,
13'b1001100000011,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1010100010011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100: edge_mask_reg_512p1[465] <= 1'b1;
 		default: edge_mask_reg_512p1[465] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000101,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110100,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110100,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b111011110100,
13'b111011110101,
13'b111011111001,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101100100,
13'b111101101001,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101100011,
13'b1000101100100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1010100010011,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100: edge_mask_reg_512p1[466] <= 1'b1;
 		default: edge_mask_reg_512p1[466] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010110,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100110,
13'b1100101010,
13'b1100101011,
13'b1100110110,
13'b1100110111,
13'b1100111010,
13'b1100111011,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100101,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100100,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100100,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b110011101001,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b110110001010,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101011001,
13'b111101011010,
13'b111101100011,
13'b111101101001,
13'b111101101010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110011,
13'b1000100110100,
13'b1000101000011,
13'b1000101000100,
13'b1000101010011,
13'b1000101010100,
13'b1000101100011,
13'b1001100110011,
13'b1001101000011,
13'b1001101010011: edge_mask_reg_512p1[467] <= 1'b1;
 		default: edge_mask_reg_512p1[467] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010110,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100110,
13'b1100101010,
13'b1100101011,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100101,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100100,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100100,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b101011011001,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111001,
13'b110101111010,
13'b110110001010,
13'b111011111001,
13'b111011111010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101010011,
13'b111101010100,
13'b111101011001,
13'b111101011010,
13'b111101100011,
13'b111101101001,
13'b111101101010,
13'b1000100000100,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101010011,
13'b1000101010100,
13'b1000101100011,
13'b1001100010011,
13'b1001100100011,
13'b1001100110011,
13'b1001100110100,
13'b1001101000011,
13'b1001101010011: edge_mask_reg_512p1[468] <= 1'b1;
 		default: edge_mask_reg_512p1[468] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011111010,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1011011010100,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100: edge_mask_reg_512p1[469] <= 1'b1;
 		default: edge_mask_reg_512p1[469] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b111010010100,
13'b111010010101,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000100,
13'b1001100000101,
13'b1001100010100,
13'b1001100010101,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1011010110100,
13'b1011011000100,
13'b1011011010100,
13'b1011011100100,
13'b1011011110100: edge_mask_reg_512p1[470] <= 1'b1;
 		default: edge_mask_reg_512p1[470] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000100,
13'b1001100000101,
13'b1001100010100,
13'b1001100010101,
13'b1010010100011,
13'b1010010100100,
13'b1010010110011,
13'b1010010110100,
13'b1010011000011,
13'b1010011000100,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1011010110100,
13'b1011011000100,
13'b1011011010100,
13'b1011011100100,
13'b1011011110100: edge_mask_reg_512p1[471] <= 1'b1;
 		default: edge_mask_reg_512p1[471] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100100,
13'b1000100100101,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1011011010100,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[472] <= 1'b1;
 		default: edge_mask_reg_512p1[472] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1011011010100,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[473] <= 1'b1;
 		default: edge_mask_reg_512p1[473] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100101,
13'b1000100100110,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100101,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100010100,
13'b1011011010100,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[474] <= 1'b1;
 		default: edge_mask_reg_512p1[474] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100101,
13'b1000100100110,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100100101,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011011010100,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[475] <= 1'b1;
 		default: edge_mask_reg_512p1[475] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100101,
13'b1000100100110,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011011010100,
13'b1011011100100,
13'b1011011110100,
13'b1011100000100,
13'b1011100010100: edge_mask_reg_512p1[476] <= 1'b1;
 		default: edge_mask_reg_512p1[476] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100101,
13'b1000100100110,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011011010100,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101: edge_mask_reg_512p1[477] <= 1'b1;
 		default: edge_mask_reg_512p1[477] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100101,
13'b1000100100110,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010011,
13'b1010011010100,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1010100010101,
13'b1011011010100,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1100011100100,
13'b1100011110100,
13'b1100100000100: edge_mask_reg_512p1[478] <= 1'b1;
 		default: edge_mask_reg_512p1[478] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010111001,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111001,
13'b110011111010,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011011001,
13'b111011011010,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1011010000100,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1011010110101,
13'b1011011000100,
13'b1100010010100,
13'b1100010010101,
13'b1100010100100,
13'b1100010100101,
13'b1100010110100,
13'b1100010110101,
13'b1101010010101: edge_mask_reg_512p1[479] <= 1'b1;
 		default: edge_mask_reg_512p1[479] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011010,
13'b1010101010,
13'b1010111001,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001010,
13'b1100001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010011001,
13'b10010011010,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111001,
13'b11011111010,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111001,
13'b100011111010,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b111001110101,
13'b111001110110,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011001,
13'b111010011010,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000101,
13'b1001011000110,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000101,
13'b1010011000110,
13'b1011010000100,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110100,
13'b1011010110101,
13'b1100010010100,
13'b1100010010101,
13'b1100010100100,
13'b1100010100101,
13'b1100010110100,
13'b1100010110101,
13'b1101010010101: edge_mask_reg_512p1[480] <= 1'b1;
 		default: edge_mask_reg_512p1[480] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000101,
13'b110110000110,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110000101,
13'b111110000110,
13'b111110001001,
13'b111110001010,
13'b111110011001,
13'b111110011010,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000101,
13'b1001110000110,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1011100100100,
13'b1011100100101,
13'b1011100110100,
13'b1011100110101,
13'b1011101000100,
13'b1011101000101,
13'b1011101010100,
13'b1011101010101,
13'b1011101100100,
13'b1011101100101,
13'b1011101110100,
13'b1100100110101,
13'b1100101000100,
13'b1100101000101,
13'b1100101010100,
13'b1100101010101,
13'b1100101100100: edge_mask_reg_512p1[481] <= 1'b1;
 		default: edge_mask_reg_512p1[481] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b101010111001,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1011100010100,
13'b1011100100100: edge_mask_reg_512p1[482] <= 1'b1;
 		default: edge_mask_reg_512p1[482] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011101001,
13'b111011101010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b111101001010,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1011100010100,
13'b1011100100100: edge_mask_reg_512p1[483] <= 1'b1;
 		default: edge_mask_reg_512p1[483] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b101010101001,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b111011000100,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b1000011010011,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1011100000100,
13'b1011100010100,
13'b1011100100100: edge_mask_reg_512p1[484] <= 1'b1;
 		default: edge_mask_reg_512p1[484] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b111011000100,
13'b111011000101,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011011001,
13'b111011011010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101001001,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1001011100011,
13'b1001011100100,
13'b1001011110011,
13'b1001011110100,
13'b1001100000011,
13'b1001100000100,
13'b1001100010011,
13'b1001100010100,
13'b1001100100011,
13'b1001100100100,
13'b1001100110011,
13'b1001100110100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110011,
13'b1010011110100,
13'b1010100000011,
13'b1010100000100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1011100000100,
13'b1011100010100,
13'b1011100100100: edge_mask_reg_512p1[485] <= 1'b1;
 		default: edge_mask_reg_512p1[485] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101011,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011010,
13'b11100011011,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010101100,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011001100,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011011100,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011010,
13'b111010001010,
13'b111010001011,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101000,
13'b111011101010,
13'b111011101011,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b1000010010111,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011011010,
13'b1000011101000,
13'b1001010100110,
13'b1001010100111,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100111,
13'b1001011101000,
13'b1010010100110,
13'b1010010100111,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100110,
13'b1010011100111,
13'b1011010100110,
13'b1011010100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100110,
13'b1011011100111,
13'b1100010110110,
13'b1100010110111,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100110,
13'b1101011000110,
13'b1101011000111,
13'b1101011010110,
13'b1101011010111,
13'b1101011100110,
13'b1110011000110,
13'b1110011010110,
13'b1110011100110: edge_mask_reg_512p1[486] <= 1'b1;
 		default: edge_mask_reg_512p1[486] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011010,
13'b11100011011,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011010,
13'b101100011011,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010101100,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011001100,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011011100,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b111010001010,
13'b111010001011,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101000,
13'b111011101010,
13'b111011101011,
13'b111011111010,
13'b111011111011,
13'b1000010010111,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011101000,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011101000,
13'b1010010100110,
13'b1010010100111,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100110,
13'b1011010100110,
13'b1011010100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100110,
13'b1100010110110,
13'b1100010110111,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100110,
13'b1101010110110,
13'b1101011000110,
13'b1101011000111,
13'b1101011010110,
13'b1101011010111,
13'b1101011100110,
13'b1110011000110,
13'b1110011010110: edge_mask_reg_512p1[487] <= 1'b1;
 		default: edge_mask_reg_512p1[487] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101010,
13'b1010101011,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b11001011001,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011010,
13'b11100011011,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100001111100,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011010,
13'b100100011011,
13'b101001001010,
13'b101001011010,
13'b101001011011,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101001111100,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010001100,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011010,
13'b101100011011,
13'b110001011010,
13'b110001011011,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010001100,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010011100,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010101100,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110010111100,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011001100,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011011100,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001010,
13'b110100001011,
13'b111001101010,
13'b111001101011,
13'b111001111010,
13'b111001111011,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101010,
13'b111011101011,
13'b111011111010,
13'b111011111011,
13'b1000001111000,
13'b1000010000111,
13'b1000010001000,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010011010,
13'b1000010011011,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010101010,
13'b1000010101011,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1001010000111,
13'b1001010001000,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1010010000110,
13'b1010010000111,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100110,
13'b1011010000111,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100110,
13'b1100010010110,
13'b1100010010111,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011100110,
13'b1101010100110,
13'b1101010110110,
13'b1101010110111,
13'b1101011000110,
13'b1101011000111,
13'b1101011010110,
13'b1101011100110: edge_mask_reg_512p1[488] <= 1'b1;
 		default: edge_mask_reg_512p1[488] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1100011010100,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000100,
13'b1100100000101: edge_mask_reg_512p1[489] <= 1'b1;
 		default: edge_mask_reg_512p1[489] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101011001,
13'b100101011010,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1100011010100,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000100,
13'b1100100000101: edge_mask_reg_512p1[490] <= 1'b1;
 		default: edge_mask_reg_512p1[490] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1100011010100,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000100,
13'b1100100000101: edge_mask_reg_512p1[491] <= 1'b1;
 		default: edge_mask_reg_512p1[491] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1011100010101,
13'b1100011010100,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000100,
13'b1100100000101: edge_mask_reg_512p1[492] <= 1'b1;
 		default: edge_mask_reg_512p1[492] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1100011010100,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000100,
13'b1100100000101: edge_mask_reg_512p1[493] <= 1'b1;
 		default: edge_mask_reg_512p1[493] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100101,
13'b1010100100110,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1100011010100,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000100,
13'b1100100000101: edge_mask_reg_512p1[494] <= 1'b1;
 		default: edge_mask_reg_512p1[494] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100101,
13'b1010100100110,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1100011010100,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000101: edge_mask_reg_512p1[495] <= 1'b1;
 		default: edge_mask_reg_512p1[495] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100111,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010101,
13'b1001100010110,
13'b1001100100101,
13'b1001100100110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100100101,
13'b1010100100110,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010100,
13'b1100011010100,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000101: edge_mask_reg_512p1[496] <= 1'b1;
 		default: edge_mask_reg_512p1[496] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b10101011011,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100110,
13'b110100100111,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001001,
13'b111011001010,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100111001,
13'b111100111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1001011000101,
13'b1001011000110,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010101,
13'b1010100010110,
13'b1010100100101,
13'b1010100100110,
13'b1011011010100,
13'b1011011010101,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1100011010100,
13'b1100011010101,
13'b1100011100100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100100000101: edge_mask_reg_512p1[497] <= 1'b1;
 		default: edge_mask_reg_512p1[497] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b111101111001,
13'b111101111010,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100100,
13'b1010101100101,
13'b1011100010110,
13'b1011100010111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101100100,
13'b1011101100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1100101100101,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010101,
13'b1101101010110,
13'b1110100110110: edge_mask_reg_512p1[498] <= 1'b1;
 		default: edge_mask_reg_512p1[498] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011011,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001010,
13'b10101001011,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b111100101010,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001010,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000111,
13'b1000100001000,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000110,
13'b1001100000111,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010101,
13'b1011100010110,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000101,
13'b1100100000110,
13'b1100100010101,
13'b1100100010110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100101,
13'b1101011100110,
13'b1101011110101,
13'b1101011110110,
13'b1101100000101,
13'b1101100000110,
13'b1110011010110,
13'b1110011100110: edge_mask_reg_512p1[499] <= 1'b1;
 		default: edge_mask_reg_512p1[499] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010110000100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[500] <= 1'b1;
 		default: edge_mask_reg_512p1[500] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101001,
13'b100110101010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101001,
13'b110110101010,
13'b111100001001,
13'b111100001010,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111001,
13'b111100111010,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101001010,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011001,
13'b111101011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101001,
13'b111101101010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111101111010,
13'b111110001001,
13'b111110001010,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110100,
13'b1010101110101,
13'b1010110000100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100,
13'b1011101100100,
13'b1011101110100: edge_mask_reg_512p1[501] <= 1'b1;
 		default: edge_mask_reg_512p1[501] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011010,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001010,
13'b10101001011,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101011111100,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111001,
13'b101100111010,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110101,
13'b110010110110,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011001100,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011011100,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011101100,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110011111100,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b111010101001,
13'b111010101010,
13'b111010110101,
13'b111010110110,
13'b111010111001,
13'b111010111010,
13'b111011000101,
13'b111011000110,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100000100,
13'b111100000101,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010100,
13'b111100010101,
13'b111100011001,
13'b111100011010,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011011010,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011101010,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1001011000101,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001100000100,
13'b1001100000101,
13'b1001100010100,
13'b1010011010100,
13'b1010011100100,
13'b1010011100101,
13'b1010011110100,
13'b1010011110101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010100,
13'b1011011100100,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011100000100: edge_mask_reg_512p1[502] <= 1'b1;
 		default: edge_mask_reg_512p1[502] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b10001101000,
13'b10001101001,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101001,
13'b101010101010,
13'b101010111001,
13'b101010111010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001001011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001011011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001101011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010010101,
13'b110010011001,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b111000101001,
13'b111000110101,
13'b111000110110,
13'b111000111001,
13'b111000111010,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001001010,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011001,
13'b111001011010,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101001,
13'b111001101010,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111001,
13'b111001111010,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001001,
13'b111010001010,
13'b111010010101,
13'b111010011001,
13'b111010011010,
13'b1000000100110,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000101,
13'b1000010000110,
13'b1000010010101,
13'b1001000100101,
13'b1001000110100,
13'b1001000110101,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110100,
13'b1001001110101,
13'b1001010000101,
13'b1010000110100,
13'b1010000110101,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001010100,
13'b1010001010101,
13'b1010001100100,
13'b1010001100101,
13'b1010001110100,
13'b1010001110101,
13'b1011000100100,
13'b1011000110100,
13'b1011001000100,
13'b1011001010100,
13'b1011001100100,
13'b1011001110100: edge_mask_reg_512p1[503] <= 1'b1;
 		default: edge_mask_reg_512p1[503] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001101001,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101011,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101010,
13'b101001101010,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010011100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b111010001010,
13'b111010001011,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100001010,
13'b1000010011000,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011101000,
13'b1000011101001,
13'b1001010011000,
13'b1001010100111,
13'b1001010101000,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011101000,
13'b1010010010111,
13'b1010010011000,
13'b1010010100111,
13'b1010010101000,
13'b1010010110111,
13'b1010010111000,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1010011100111,
13'b1010011101000,
13'b1011010010111,
13'b1011010100111,
13'b1011010101000,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010111,
13'b1011011011000,
13'b1011011100111,
13'b1011011101000,
13'b1100010010111,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1101010100111,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1101011100110,
13'b1101011100111,
13'b1101011101000,
13'b1110010110110,
13'b1110010110111,
13'b1110011000110,
13'b1110011000111,
13'b1110011010110,
13'b1110011010111,
13'b1110011100110,
13'b1110011100111,
13'b1111010110110,
13'b1111011000110,
13'b1111011000111,
13'b1111011010110,
13'b1111011010111,
13'b1111011100110,
13'b1111011100111: edge_mask_reg_512p1[504] <= 1'b1;
 		default: edge_mask_reg_512p1[504] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001011,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b101001111010,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b1000010100111,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001010,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011010,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110111,
13'b1000011111000,
13'b1001010100110,
13'b1001010100111,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110111,
13'b1001011111000,
13'b1010010100110,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110110,
13'b1010011110111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110110,
13'b1011011110111,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1101011000110,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011100101,
13'b1101011100110,
13'b1101011100111,
13'b1101011110101,
13'b1101011110110,
13'b1101100000110,
13'b1110011010101,
13'b1110011010110,
13'b1110011100101,
13'b1110011100110,
13'b1110011110110,
13'b1110100000110,
13'b1111011100110,
13'b1111011110110: edge_mask_reg_512p1[505] <= 1'b1;
 		default: edge_mask_reg_512p1[505] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001011,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b1000010100110,
13'b1000010100111,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011010,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110111,
13'b1000011111000,
13'b1001010100110,
13'b1001010100111,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110111,
13'b1001011111000,
13'b1010010100110,
13'b1010010100111,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110110,
13'b1010011110111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011100110,
13'b1011011100111,
13'b1011011110110,
13'b1011011110111,
13'b1100010110110,
13'b1100010110111,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1101011000110,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011100101,
13'b1101011100110,
13'b1101011100111,
13'b1101011110101,
13'b1101011110110,
13'b1101100000110,
13'b1110011010110,
13'b1110011100101,
13'b1110011100110,
13'b1110011110110,
13'b1110100000110,
13'b1111011100110,
13'b1111011110110: edge_mask_reg_512p1[506] <= 1'b1;
 		default: edge_mask_reg_512p1[506] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111001,
13'b10111010,
13'b11001001,
13'b11001010,
13'b11011001,
13'b11011010,
13'b11101001,
13'b11101010,
13'b11111001,
13'b11111010,
13'b100001001,
13'b100001010,
13'b100011001,
13'b100011010,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111001,
13'b1010001001,
13'b1010001010,
13'b1010011001,
13'b1010011010,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111011,
13'b10001101001,
13'b10001111001,
13'b10001111010,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101011,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101010,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010101100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b111010001001,
13'b111010001010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100001010,
13'b1000010100111,
13'b1000010101000,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011101000,
13'b1000011101001,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011101000,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010111,
13'b1010011011000,
13'b1010011100111,
13'b1010011101000,
13'b1011010100110,
13'b1011010100111,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100111,
13'b1011011101000,
13'b1100010100111,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1101010110110,
13'b1101010110111,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1101011100110,
13'b1101011100111,
13'b1101011101000,
13'b1110011000110,
13'b1110011000111,
13'b1110011010110,
13'b1110011010111,
13'b1110011100110,
13'b1110011100111,
13'b1111011000110,
13'b1111011010110,
13'b1111011010111,
13'b1111011100110,
13'b1111011100111: edge_mask_reg_512p1[507] <= 1'b1;
 		default: edge_mask_reg_512p1[507] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111011,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101011,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101010,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001010,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100111,
13'b1000011101000,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100101,
13'b1101011100110,
13'b1101011110101,
13'b1101011110110,
13'b1110011010101,
13'b1110011010110,
13'b1110011100101,
13'b1110011100110: edge_mask_reg_512p1[508] <= 1'b1;
 		default: edge_mask_reg_512p1[508] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111011,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001111010,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101010111100,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011001100,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011011100,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011101100,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010101011,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b1000010100111,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001010,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011010,
13'b1000011100111,
13'b1000011101000,
13'b1001010100110,
13'b1001010100111,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1010010100110,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1011010110110,
13'b1011010110111,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1101011000101,
13'b1101011000110,
13'b1101011010101,
13'b1101011010110,
13'b1101011100101,
13'b1101011100110,
13'b1101011110101,
13'b1101011110110,
13'b1110011010101,
13'b1110011010110,
13'b1110011100101,
13'b1110011100110: edge_mask_reg_512p1[509] <= 1'b1;
 		default: edge_mask_reg_512p1[509] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b101001010,
13'b1001111000,
13'b1001111001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011010,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001011,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b110010001001,
13'b110010001010,
13'b110010011001,
13'b110010011010,
13'b110010101001,
13'b110010101010,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b111010011001,
13'b111010011010,
13'b111010101001,
13'b111010101010,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100001001,
13'b111100001010,
13'b111100011001,
13'b111100011010,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110111,
13'b1000011111000,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110111,
13'b1001011111000,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110110,
13'b1010011110111,
13'b1011010110110,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110110,
13'b1011011110111,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011100101,
13'b1101011100110,
13'b1101011100111,
13'b1101011110101,
13'b1101011110110,
13'b1101100000110,
13'b1110011010101,
13'b1110011010110,
13'b1110011100101,
13'b1110011100110,
13'b1110011110110,
13'b1110100000110,
13'b1111011100110,
13'b1111011110110: edge_mask_reg_512p1[510] <= 1'b1;
 		default: edge_mask_reg_512p1[510] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101001,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110100,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b110011011001,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110100,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001001,
13'b111011101001,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111001,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100001001,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101001000,
13'b111101001001,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101011001,
13'b111101100100,
13'b111101101001,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101100011,
13'b1000101100100,
13'b1001011110100,
13'b1001011110101,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101010011,
13'b1001101010100,
13'b1001101100011,
13'b1001101100100,
13'b1010100010011,
13'b1010100010100,
13'b1010100100011,
13'b1010100100100,
13'b1010100110011,
13'b1010100110100,
13'b1010101000011,
13'b1010101000100,
13'b1010101010011,
13'b1010101010100,
13'b1010101100011,
13'b1010101100100,
13'b1011100010100,
13'b1011100100100,
13'b1011100110100,
13'b1011101000100,
13'b1011101010100,
13'b1100100100100: edge_mask_reg_512p1[511] <= 1'b1;
 		default: edge_mask_reg_512p1[511] <= 1'b0;
 	endcase

end
endmodule

