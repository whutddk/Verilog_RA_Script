/*******************************************
****** Wuhan university of technology ******
****** Ruige Lee ******
year: 2019
month: 3
date: 4
hour: 17
minutes: 7
second: 2
********************************************/

module prm_LUTX1_Sp_3_4_4_chk512p7(
	input [2:0] x,
	input [3:0] y,
	input [3:0] z,
	output [511:0] edge_mask_512p7
);

	reg [511:0] edge_mask_reg_512p7;
	assign edge_mask_512p7= edge_mask_reg_512p7;

always @( *) begin
    case({x,y,z})
		default: edge_mask_reg_512p7[0] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[1] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[2] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[3] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[4] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010100111,
11'b10010101000,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011101000,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111101000,
11'b11010100110,
11'b11010100111,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010111,
11'b11011011000,
11'b11011101000,
11'b11110100110,
11'b11110100111,
11'b11110110110,
11'b11110110111,
11'b11110111000,
11'b11111000110,
11'b11111000111,
11'b11111001000,
11'b11111010111,
11'b11111011000,
11'b11111101000: edge_mask_reg_512p7[5] <= 1'b1;
 		default: edge_mask_reg_512p7[5] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[6] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111010,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001010,
11'b110001011,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111001,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010101,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110110,
11'b10011110111,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111110101,
11'b10111110110,
11'b11010100101,
11'b11010100110,
11'b11010110101,
11'b11010110110,
11'b11011000101,
11'b11011000110,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11111010101: edge_mask_reg_512p7[7] <= 1'b1;
 		default: edge_mask_reg_512p7[7] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b1000111100,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111011,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001101100,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010011001,
11'b10101011001,
11'b10101101001,
11'b10101101010,
11'b10101111000,
11'b10101111001,
11'b10101111010,
11'b10110001000,
11'b10110001001,
11'b10110001010,
11'b10110011000,
11'b10110011001,
11'b11001101000,
11'b11001101001,
11'b11001101010,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11001111010,
11'b11010000111,
11'b11010001000,
11'b11010001001,
11'b11010011000,
11'b11010011001,
11'b11101101000,
11'b11101101001,
11'b11101110111,
11'b11101111000,
11'b11101111001,
11'b11110000111,
11'b11110001000,
11'b11110001001: edge_mask_reg_512p7[8] <= 1'b1;
 		default: edge_mask_reg_512p7[8] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1101000101,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010100,
11'b1110010101,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101010,
11'b10001000101,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111010,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001010,
11'b10010010100,
11'b10010010101,
11'b10101100101,
11'b10101100110,
11'b10101110100,
11'b10101110101,
11'b10101110110: edge_mask_reg_512p7[9] <= 1'b1;
 		default: edge_mask_reg_512p7[9] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100111000,
11'b1100111001,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100110,
11'b10100000110,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b11000000101,
11'b11000000110,
11'b11000010100,
11'b11000010101,
11'b11000010110,
11'b11000100100,
11'b11000100101,
11'b11000100110,
11'b11100010100,
11'b11100010101: edge_mask_reg_512p7[10] <= 1'b1;
 		default: edge_mask_reg_512p7[10] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[11] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101011,
11'b101111011,
11'b101111100,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b111001011,
11'b1001111100,
11'b1001111101,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001011,
11'b1011001100,
11'b1011011011,
11'b1011011100,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b1111011011,
11'b1111011100,
11'b10010101011,
11'b10010101100,
11'b10010111011,
11'b10010111100,
11'b10011001011,
11'b10011001100,
11'b10011011011,
11'b10011011100,
11'b10110101011,
11'b10110101100,
11'b10110111011,
11'b10110111100,
11'b10111001011,
11'b10111001100,
11'b10111011011,
11'b10111011100,
11'b11010101011,
11'b11010111010,
11'b11010111011,
11'b11010111100,
11'b11011001010,
11'b11011001011,
11'b11011001100,
11'b11011011011,
11'b11011011100,
11'b11110101010,
11'b11110101011,
11'b11110111010,
11'b11110111011,
11'b11111001010,
11'b11111001011,
11'b11111011010,
11'b11111011011: edge_mask_reg_512p7[12] <= 1'b1;
 		default: edge_mask_reg_512p7[12] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[13] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001011,
11'b1000011000,
11'b1000011001,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1100010101,
11'b1100010110,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b10000010100,
11'b10000100100,
11'b10000100101,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10001000100,
11'b10001000101,
11'b10001001010,
11'b10001010100,
11'b10001010101,
11'b10001011010,
11'b10100100011,
11'b10100100100,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10101000100,
11'b10101000101,
11'b10101010100,
11'b10101010101: edge_mask_reg_512p7[14] <= 1'b1;
 		default: edge_mask_reg_512p7[14] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111001,
11'b10111010,
11'b11001000,
11'b11001001,
11'b11001010,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111001001,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111001,
11'b10011010101,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10011110101,
11'b10011110110,
11'b10011110111,
11'b10111100100,
11'b10111100101,
11'b10111100110,
11'b10111110100,
11'b10111110101,
11'b10111110110,
11'b11011100100,
11'b11011110100: edge_mask_reg_512p7[15] <= 1'b1;
 		default: edge_mask_reg_512p7[15] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010101010,
11'b1010101011,
11'b1010110110,
11'b1010110111,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110101010,
11'b1110101011,
11'b1110110101,
11'b1110110110,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111001,
11'b10011000101,
11'b10011000110,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011010111,
11'b10011011010,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10011101010,
11'b10011110101,
11'b10011110110,
11'b10011110111,
11'b10111010100,
11'b10111010101,
11'b10111100100,
11'b10111100101,
11'b10111100110,
11'b10111110100,
11'b10111110101,
11'b10111110110: edge_mask_reg_512p7[16] <= 1'b1;
 		default: edge_mask_reg_512p7[16] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111011,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010100,
11'b1111010101,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111001,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011101010,
11'b10011110101,
11'b10011110110,
11'b10011111010: edge_mask_reg_512p7[17] <= 1'b1;
 		default: edge_mask_reg_512p7[17] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[18] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[19] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111001001,
11'b1111001010,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111111000,
11'b1111111001,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011111000,
11'b10011111001,
11'b10011111010,
11'b10111011000,
11'b10111011001,
11'b10111101000,
11'b10111101001,
11'b10111111000,
11'b10111111001,
11'b11011011000,
11'b11011011001,
11'b11011101000,
11'b11011101001,
11'b11011111000,
11'b11011111001,
11'b11111011000,
11'b11111011001,
11'b11111101000,
11'b11111101001,
11'b11111111000,
11'b11111111001: edge_mask_reg_512p7[20] <= 1'b1;
 		default: edge_mask_reg_512p7[20] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001010,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110100,
11'b110110101,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111001,
11'b1110111010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001111010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010001010: edge_mask_reg_512p7[21] <= 1'b1;
 		default: edge_mask_reg_512p7[21] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[22] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[23] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b1000010111,
11'b1000011000,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110110,
11'b1001110111,
11'b1100010111,
11'b1100011000,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b10000100111,
11'b10000101000,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010110,
11'b10001010111,
11'b10100100111,
11'b10100101000,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010110,
11'b10101010111,
11'b11000100111,
11'b11000101000,
11'b11000110101,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11100100110,
11'b11100100111,
11'b11100101000,
11'b11100110110,
11'b11100110111,
11'b11100111000,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101001000,
11'b11101010101,
11'b11101010110,
11'b11101010111: edge_mask_reg_512p7[24] <= 1'b1;
 		default: edge_mask_reg_512p7[24] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b10000010111,
11'b10000011000,
11'b10000100111,
11'b10000101000,
11'b10000110111,
11'b10000111000,
11'b10100000111,
11'b10100001000,
11'b10100010111,
11'b10100011000,
11'b10100100111,
11'b10100101000,
11'b10100110111,
11'b10100111000,
11'b11000000111,
11'b11000010110,
11'b11000010111,
11'b11000011000,
11'b11000100110,
11'b11000100111,
11'b11000101000,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11100000111,
11'b11100010110,
11'b11100010111,
11'b11100011000,
11'b11100100110,
11'b11100100111,
11'b11100101000,
11'b11100110110,
11'b11100110111,
11'b11100111000: edge_mask_reg_512p7[25] <= 1'b1;
 		default: edge_mask_reg_512p7[25] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10001010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101101000,
11'b1101101001,
11'b10000011000,
11'b10000100111,
11'b10000101000,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10001001000,
11'b10001001001,
11'b10001011000,
11'b10001011001,
11'b10100010111,
11'b10100011000,
11'b10100100111,
11'b10100101000,
11'b10100110111,
11'b10100111000,
11'b10101000111,
11'b10101001000,
11'b10101001001,
11'b10101011000,
11'b10101011001,
11'b11000010111,
11'b11000011000,
11'b11000100110,
11'b11000100111,
11'b11000101000,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001001001,
11'b11001010111,
11'b11001011000,
11'b11001011001,
11'b11100010111,
11'b11100100110,
11'b11100100111,
11'b11100101000,
11'b11100110110,
11'b11100110111,
11'b11100111000,
11'b11101000110,
11'b11101000111,
11'b11101001000,
11'b11101001001,
11'b11101010111,
11'b11101011000,
11'b11101011001: edge_mask_reg_512p7[26] <= 1'b1;
 		default: edge_mask_reg_512p7[26] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100111,
11'b1101101000,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10100010100,
11'b10100010101,
11'b10100100100,
11'b10100100101,
11'b10100110100,
11'b10100110101,
11'b10101000100,
11'b10101000101,
11'b10101010100,
11'b10101010101,
11'b11000010100,
11'b11000010101,
11'b11000100100,
11'b11000100101,
11'b11000110100,
11'b11000110101,
11'b11001000100,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11100100100,
11'b11100110100,
11'b11101000100: edge_mask_reg_512p7[27] <= 1'b1;
 		default: edge_mask_reg_512p7[27] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100011,
11'b10001100100,
11'b10100010100,
11'b10100010101,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101100011,
11'b11000010100,
11'b11000010101,
11'b11000100100,
11'b11000100101,
11'b11000110100,
11'b11000110101: edge_mask_reg_512p7[28] <= 1'b1;
 		default: edge_mask_reg_512p7[28] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10100010100,
11'b10100010101,
11'b10100100100,
11'b10100100101,
11'b10100110100,
11'b10100110101,
11'b11000000101,
11'b11000010100,
11'b11000010101,
11'b11000100100,
11'b11000100101,
11'b11000110100,
11'b11000110101,
11'b11100010100,
11'b11100100100: edge_mask_reg_512p7[29] <= 1'b1;
 		default: edge_mask_reg_512p7[29] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101101000,
11'b1101101001,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010110,
11'b10001010111,
11'b10100010100,
11'b10100010101,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b10101010110,
11'b11000010100,
11'b11000010101,
11'b11000100100,
11'b11000100101,
11'b11000100110,
11'b11000110100,
11'b11000110101,
11'b11000110110,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010101,
11'b11001010110,
11'b11100100100,
11'b11100100101,
11'b11100110100,
11'b11100110101,
11'b11100110110,
11'b11101000100,
11'b11101000101,
11'b11101000110: edge_mask_reg_512p7[30] <= 1'b1;
 		default: edge_mask_reg_512p7[30] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001010,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110101001,
11'b1110101010,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10110110110,
11'b10110110111,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b11011000101,
11'b11011000110,
11'b11011000111,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11111000101,
11'b11111000110,
11'b11111010101,
11'b11111010110,
11'b11111100101,
11'b11111100110: edge_mask_reg_512p7[31] <= 1'b1;
 		default: edge_mask_reg_512p7[31] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111000110,
11'b10111010110,
11'b10111010111,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111010101,
11'b11111010110,
11'b11111100101,
11'b11111100110,
11'b11111110101,
11'b11111110110,
11'b11111110111: edge_mask_reg_512p7[32] <= 1'b1;
 		default: edge_mask_reg_512p7[32] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10011110111,
11'b10011111000,
11'b10011111001,
11'b10111000110,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11011111000,
11'b11111010101,
11'b11111010110,
11'b11111100101,
11'b11111100110,
11'b11111100111,
11'b11111110110,
11'b11111110111: edge_mask_reg_512p7[33] <= 1'b1;
 		default: edge_mask_reg_512p7[33] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010011011,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110101010,
11'b1110101011,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10010111000,
11'b10010111001,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10110111000,
11'b10110111001,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b11010110111,
11'b11010111000,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011101000,
11'b11111000110,
11'b11111000111,
11'b11111001000,
11'b11111010101,
11'b11111010110,
11'b11111010111,
11'b11111011000,
11'b11111100101,
11'b11111100110: edge_mask_reg_512p7[34] <= 1'b1;
 		default: edge_mask_reg_512p7[34] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011100110,
11'b1011100111,
11'b11011110101,
11'b11011110110: edge_mask_reg_512p7[35] <= 1'b1;
 		default: edge_mask_reg_512p7[35] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[36] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001010,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001010,
11'b111001011,
11'b111011010,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101010,
11'b1110001011,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101010,
11'b1111101011,
11'b10010101010,
11'b10010101011,
11'b10010111001,
11'b10010111010,
11'b10010111011,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011101010,
11'b10110101010,
11'b10110101011,
11'b10110111001,
11'b10110111010,
11'b10110111011,
11'b10111001001,
11'b10111001010,
11'b10111001011,
11'b10111011001,
11'b10111011010,
11'b10111101001,
11'b10111101010,
11'b11010101010,
11'b11010101011,
11'b11010111001,
11'b11010111010,
11'b11010111011,
11'b11011001001,
11'b11011001010,
11'b11011011001,
11'b11011011010,
11'b11011101001,
11'b11110101010,
11'b11110111001,
11'b11110111010,
11'b11111001000,
11'b11111001001,
11'b11111001010,
11'b11111011000,
11'b11111011001,
11'b11111011010,
11'b11111101001: edge_mask_reg_512p7[37] <= 1'b1;
 		default: edge_mask_reg_512p7[37] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10100010101,
11'b10100010110: edge_mask_reg_512p7[38] <= 1'b1;
 		default: edge_mask_reg_512p7[38] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100111010,
11'b100111011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000101010,
11'b1000101011,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011011,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b10000010101,
11'b10000010110,
11'b10000010111: edge_mask_reg_512p7[39] <= 1'b1;
 		default: edge_mask_reg_512p7[39] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[40] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[41] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[42] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1000110111,
11'b1000111000,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b10001000100,
11'b10001000101,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100011,
11'b10101000100,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100011,
11'b11001010100,
11'b11001100100,
11'b11001100101,
11'b11001110100,
11'b11001110101: edge_mask_reg_512p7[43] <= 1'b1;
 		default: edge_mask_reg_512p7[43] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1000110111,
11'b1000111000,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110100111,
11'b1110101000,
11'b10001000100,
11'b10001000101,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101000100,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b10110010011,
11'b10110010100,
11'b11001010100,
11'b11001100100,
11'b11001100101,
11'b11001110100,
11'b11001110101: edge_mask_reg_512p7[44] <= 1'b1;
 		default: edge_mask_reg_512p7[44] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001010,
11'b111001011,
11'b111011010,
11'b1010011100,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101001,
11'b1011101010,
11'b1110101011,
11'b1110101100,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111111000,
11'b1111111001,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011001100,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011011100,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101011,
11'b10011111000,
11'b10011111001,
11'b10011111010,
11'b10111001000,
11'b10111001001,
11'b10111001010,
11'b10111011000,
11'b10111011001,
11'b10111011010,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b10111110111,
11'b10111111000,
11'b10111111001,
11'b11011001000,
11'b11011001001,
11'b11011001010,
11'b11011010111,
11'b11011011000,
11'b11011011001,
11'b11011100111,
11'b11011101000,
11'b11011101001,
11'b11011110111,
11'b11011111000,
11'b11111001000,
11'b11111001001,
11'b11111010111,
11'b11111011000,
11'b11111011001,
11'b11111100111,
11'b11111101000: edge_mask_reg_512p7[45] <= 1'b1;
 		default: edge_mask_reg_512p7[45] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001011,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111111001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011100111,
11'b10011101000,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100110,
11'b11011100111,
11'b11110110110,
11'b11110110111,
11'b11111000110,
11'b11111000111,
11'b11111001000,
11'b11111010110,
11'b11111010111,
11'b11111100110,
11'b11111100111: edge_mask_reg_512p7[46] <= 1'b1;
 		default: edge_mask_reg_512p7[46] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111000111,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b11011000111,
11'b11011010110,
11'b11011010111,
11'b11011100110,
11'b11011100111,
11'b11011110110,
11'b11011110111,
11'b11111010110,
11'b11111010111,
11'b11111100110,
11'b11111100111,
11'b11111110110,
11'b11111110111: edge_mask_reg_512p7[47] <= 1'b1;
 		default: edge_mask_reg_512p7[47] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111000111,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b11011000111,
11'b11011010110,
11'b11011010111,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111010110,
11'b11111010111,
11'b11111100101,
11'b11111100110,
11'b11111100111,
11'b11111110101,
11'b11111110110: edge_mask_reg_512p7[48] <= 1'b1;
 		default: edge_mask_reg_512p7[48] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111000111,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b11011000111,
11'b11011010110,
11'b11011010111,
11'b11011100110,
11'b11011100111,
11'b11011110110,
11'b11011110111,
11'b11111010110,
11'b11111010111,
11'b11111100101,
11'b11111100110,
11'b11111100111,
11'b11111110101,
11'b11111110110,
11'b11111110111: edge_mask_reg_512p7[49] <= 1'b1;
 		default: edge_mask_reg_512p7[49] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110001001,
11'b1110001010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111111001,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100111,
11'b10011101000,
11'b10110010101,
11'b10110010110,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11011000101,
11'b11011000110,
11'b11011000111,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011100110,
11'b11011100111,
11'b11110100101,
11'b11110110101,
11'b11110110110,
11'b11111000101,
11'b11111000110,
11'b11111010101,
11'b11111010110,
11'b11111010111,
11'b11111100110,
11'b11111100111: edge_mask_reg_512p7[50] <= 1'b1;
 		default: edge_mask_reg_512p7[50] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111100,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101011,
11'b1101101100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011011,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000101011,
11'b10000101100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10000111011,
11'b10000111100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10100010110,
11'b10100100110: edge_mask_reg_512p7[51] <= 1'b1;
 		default: edge_mask_reg_512p7[51] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001010,
11'b1001001011,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011011,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100100101,
11'b10100100110: edge_mask_reg_512p7[52] <= 1'b1;
 		default: edge_mask_reg_512p7[52] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100111010,
11'b100111011,
11'b1000011000,
11'b1000011001,
11'b1000101010,
11'b1000101011,
11'b1000111011,
11'b1000111100,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011011,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111011,
11'b1100111100,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10100000110,
11'b10100000111,
11'b10100001000,
11'b10100010110: edge_mask_reg_512p7[53] <= 1'b1;
 		default: edge_mask_reg_512p7[53] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100111010,
11'b100111011,
11'b1000011000,
11'b1000011001,
11'b1000101010,
11'b1000101011,
11'b1000111011,
11'b1000111100,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111011,
11'b1100111100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10100000111,
11'b10100010110: edge_mask_reg_512p7[54] <= 1'b1;
 		default: edge_mask_reg_512p7[54] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100111010,
11'b100111011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000101010,
11'b1000101011,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011011,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10100010110: edge_mask_reg_512p7[55] <= 1'b1;
 		default: edge_mask_reg_512p7[55] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111100,
11'b1100101100,
11'b1100111100: edge_mask_reg_512p7[56] <= 1'b1;
 		default: edge_mask_reg_512p7[56] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011010,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110111,
11'b10011111000,
11'b10111000110,
11'b10111000111,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111010101,
11'b11111010110,
11'b11111100101,
11'b11111100110,
11'b11111110110: edge_mask_reg_512p7[57] <= 1'b1;
 		default: edge_mask_reg_512p7[57] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011101000,
11'b1011101001,
11'b1111101001,
11'b1111101010,
11'b1111111001,
11'b10111110111,
11'b11011110111,
11'b11111110111: edge_mask_reg_512p7[58] <= 1'b1;
 		default: edge_mask_reg_512p7[58] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[59] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111111000,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101011,
11'b10011111000,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b10111110111,
11'b10111111000,
11'b11011000101,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100110,
11'b11011100111,
11'b11011101000,
11'b11011110111,
11'b11011111000,
11'b11111000110,
11'b11111010110,
11'b11111010111,
11'b11111100110,
11'b11111100111,
11'b11111101000: edge_mask_reg_512p7[60] <= 1'b1;
 		default: edge_mask_reg_512p7[60] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1010001010,
11'b1010001011,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101001,
11'b1011101010,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111111000,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011101000,
11'b10011101001,
11'b10011101011,
11'b10011111000,
11'b10110101000,
11'b10110101001,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b10111111000,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11010110111,
11'b11010111000,
11'b11010111001,
11'b11011000111,
11'b11011001000,
11'b11011001001,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100110,
11'b11011100111,
11'b11011101000,
11'b11011110111,
11'b11011111000,
11'b11110100111,
11'b11110101000,
11'b11110110111,
11'b11110111000,
11'b11111000111,
11'b11111001000,
11'b11111010111,
11'b11111011000,
11'b11111100111,
11'b11111101000: edge_mask_reg_512p7[61] <= 1'b1;
 		default: edge_mask_reg_512p7[61] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101001,
11'b1011101010,
11'b1110101011,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111111000,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101011,
11'b10011111000,
11'b10111001000,
11'b10111001001,
11'b10111001010,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111011010,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b10111101010,
11'b10111111000,
11'b11011001000,
11'b11011001001,
11'b11011010111,
11'b11011011000,
11'b11011011001,
11'b11011100110,
11'b11011100111,
11'b11011101000,
11'b11011101001,
11'b11011110111,
11'b11011111000,
11'b11111001000,
11'b11111001001,
11'b11111010111,
11'b11111011000,
11'b11111011001,
11'b11111100111,
11'b11111101000,
11'b11111101001: edge_mask_reg_512p7[62] <= 1'b1;
 		default: edge_mask_reg_512p7[62] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111011000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b10010100100,
11'b10010100101,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10110100100,
11'b10110100101,
11'b10110110100,
11'b10110110101,
11'b10111000100,
11'b10111000101,
11'b10111000110,
11'b10111010100,
11'b10111010101,
11'b10111010110,
11'b10111100101,
11'b11010100100,
11'b11010110100,
11'b11010110101,
11'b11011000100,
11'b11011000101,
11'b11011010100,
11'b11011010101,
11'b11011100101,
11'b11110110100,
11'b11110110101,
11'b11111000100,
11'b11111000101,
11'b11111010100,
11'b11111010101,
11'b11111100101: edge_mask_reg_512p7[63] <= 1'b1;
 		default: edge_mask_reg_512p7[63] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[64] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101011,
11'b10111011,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b101111011,
11'b101111100,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b111001011,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001011,
11'b1011001100,
11'b1011011011,
11'b1011011100,
11'b1101011100,
11'b1101011101,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b1111011011,
11'b1111011100,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010001100,
11'b10010001101,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10010011101,
11'b10010101001,
11'b10010101010,
11'b10010101011,
11'b10010101100,
11'b10010101101,
11'b10010111010,
11'b10010111011,
11'b10010111100,
11'b10110001001,
11'b10110001010,
11'b10110001011,
11'b10110011000,
11'b10110011001,
11'b10110011010,
11'b10110011011,
11'b10110101001,
11'b10110101010,
11'b10110101011,
11'b10110111001,
11'b10110111010,
11'b10110111011,
11'b11010001001,
11'b11010001010,
11'b11010011000,
11'b11010011001,
11'b11010011010,
11'b11010101000,
11'b11010101001,
11'b11010101010,
11'b11010111001,
11'b11010111010,
11'b11110011000,
11'b11110011001,
11'b11110011010,
11'b11110101000,
11'b11110101001,
11'b11110101010,
11'b11110111001,
11'b11110111010: edge_mask_reg_512p7[65] <= 1'b1;
 		default: edge_mask_reg_512p7[65] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101011,
11'b10111011,
11'b101101011,
11'b101101100,
11'b101111011,
11'b101111100,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b111001011,
11'b1001101100,
11'b1001101101,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001011,
11'b1011001100,
11'b1011011011,
11'b1011011100,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b1111011011,
11'b1111011100,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10010101010,
11'b10010101011,
11'b10010101100,
11'b10010101101,
11'b10010111010,
11'b10010111011,
11'b10010111100,
11'b10010111101,
11'b10011001010,
11'b10011001011,
11'b10011001100,
11'b10011001101,
11'b10011011011,
11'b10011011100,
11'b10110011001,
11'b10110011010,
11'b10110011011,
11'b10110101001,
11'b10110101010,
11'b10110101011,
11'b10110111001,
11'b10110111010,
11'b10110111011,
11'b10110111100,
11'b10111001010,
11'b10111001011,
11'b10111001100,
11'b10111011011,
11'b10111011100,
11'b11010011001,
11'b11010011010,
11'b11010101000,
11'b11010101001,
11'b11010101010,
11'b11010101011,
11'b11010111001,
11'b11010111010,
11'b11010111011,
11'b11011001010,
11'b11011001011,
11'b11011001100,
11'b11011011010,
11'b11011011011,
11'b11011011100,
11'b11110011001,
11'b11110011010,
11'b11110101000,
11'b11110101001,
11'b11110101010,
11'b11110101011,
11'b11110111001,
11'b11110111010,
11'b11110111011,
11'b11111001001,
11'b11111001010,
11'b11111001011,
11'b11111011010,
11'b11111011011: edge_mask_reg_512p7[66] <= 1'b1;
 		default: edge_mask_reg_512p7[66] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[67] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10101110100,
11'b10101110101,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11110000100,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101: edge_mask_reg_512p7[68] <= 1'b1;
 		default: edge_mask_reg_512p7[68] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b1001010111,
11'b1001011000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101100111,
11'b1101101000,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10001100101,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10101110100,
11'b10101110101,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11110000100,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101: edge_mask_reg_512p7[69] <= 1'b1;
 		default: edge_mask_reg_512p7[69] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b10010000101,
11'b10010000110,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000110,
11'b10011000111,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10111000110,
11'b10111000111,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110101,
11'b11010110110,
11'b11011000110,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101,
11'b11110100110,
11'b11110110101,
11'b11110110110: edge_mask_reg_512p7[70] <= 1'b1;
 		default: edge_mask_reg_512p7[70] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011101000,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010000101,
11'b10010000110,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11010110101,
11'b11011000100,
11'b11011000101,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101,
11'b11110110100: edge_mask_reg_512p7[71] <= 1'b1;
 		default: edge_mask_reg_512p7[71] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010111,
11'b1011011000,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000100,
11'b1111000101,
11'b1111000111,
11'b1111001000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000011,
11'b10011000100,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10111000011,
11'b10111000100,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11010110101,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101: edge_mask_reg_512p7[72] <= 1'b1;
 		default: edge_mask_reg_512p7[72] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b10010000101,
11'b10010000110,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000101,
11'b10011000110,
11'b10011010101,
11'b10011010110,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10111000100,
11'b10111000101,
11'b10111000110,
11'b10111010100,
11'b10111010101,
11'b10111010110,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11010110101,
11'b11011000100,
11'b11011000101,
11'b11011010100,
11'b11011010101,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101,
11'b11110110100,
11'b11110110101,
11'b11111000100,
11'b11111000101,
11'b11111010100,
11'b11111010101: edge_mask_reg_512p7[73] <= 1'b1;
 		default: edge_mask_reg_512p7[73] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10001110101,
11'b10001110110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10101110101,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11110000100,
11'b11110000101,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101: edge_mask_reg_512p7[74] <= 1'b1;
 		default: edge_mask_reg_512p7[74] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010000101,
11'b10010000110,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10011000110,
11'b10011000111,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10111000110,
11'b10111000111,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11011000110,
11'b11011000111,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101,
11'b11110100110,
11'b11110110101,
11'b11110110110,
11'b11111000101,
11'b11111000110: edge_mask_reg_512p7[75] <= 1'b1;
 		default: edge_mask_reg_512p7[75] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010111,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000011,
11'b10011000100,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10111000011,
11'b10111000100,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11010110101,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101: edge_mask_reg_512p7[76] <= 1'b1;
 		default: edge_mask_reg_512p7[76] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10011001,
11'b10011010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000010111,
11'b1000011000,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110001000,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b11000100100,
11'b11000100101,
11'b11000110100,
11'b11000110101,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100101,
11'b11001100110,
11'b11100110100,
11'b11101000100,
11'b11101000101,
11'b11101010100,
11'b11101010101,
11'b11101010110,
11'b11101100101,
11'b11101100110: edge_mask_reg_512p7[77] <= 1'b1;
 		default: edge_mask_reg_512p7[77] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10011001,
11'b10011010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100111000,
11'b1100111001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110001000,
11'b1110001001,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b11001000110,
11'b11001000111,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100101,
11'b11001100110,
11'b11101000101,
11'b11101000110,
11'b11101010101,
11'b11101010110,
11'b11101100101,
11'b11101100110: edge_mask_reg_512p7[78] <= 1'b1;
 		default: edge_mask_reg_512p7[78] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110011000,
11'b1110011001,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b11001010101,
11'b11001010110,
11'b11001100101,
11'b11001100110,
11'b11001110101,
11'b11001110110,
11'b11010000101,
11'b11010000110,
11'b11101010101,
11'b11101010110,
11'b11101100101,
11'b11101100110,
11'b11101110101,
11'b11101110110,
11'b11110000101,
11'b11110000110: edge_mask_reg_512p7[79] <= 1'b1;
 		default: edge_mask_reg_512p7[79] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010111010,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10110111010,
11'b10110111011,
11'b10111001001,
11'b10111001010,
11'b10111001011,
11'b10111011010,
11'b10111011011,
11'b11010111010,
11'b11010111011,
11'b11011001010,
11'b11011001011,
11'b11011011010,
11'b11011011011,
11'b11110111010,
11'b11110111011,
11'b11111001010,
11'b11111001011,
11'b11111011010,
11'b11111011011: edge_mask_reg_512p7[80] <= 1'b1;
 		default: edge_mask_reg_512p7[80] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[81] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[82] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111010110,
11'b111010111,
11'b111011000,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011010110,
11'b1011010111,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000100,
11'b1111000110,
11'b1111000111,
11'b10010000100,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000100,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10111000011,
11'b10111000100,
11'b11010010100,
11'b11010100100,
11'b11010110100: edge_mask_reg_512p7[83] <= 1'b1;
 		default: edge_mask_reg_512p7[83] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b10010000100,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10110010011,
11'b10110010100,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111000110,
11'b10111010100,
11'b10111010101,
11'b10111010110,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11010110101,
11'b11011000100,
11'b11011000101,
11'b11011010100,
11'b11011010101,
11'b11110110100,
11'b11110110101,
11'b11111000100,
11'b11111000101,
11'b11111010100,
11'b11111010101: edge_mask_reg_512p7[84] <= 1'b1;
 		default: edge_mask_reg_512p7[84] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100101,
11'b1100110,
11'b1100111,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000110,
11'b1111000111,
11'b10010000011,
11'b10010000100,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10110000011,
11'b10110000100,
11'b10110010011,
11'b10110010100,
11'b10110100011,
11'b10110100100,
11'b10110110011,
11'b10110110100: edge_mask_reg_512p7[85] <= 1'b1;
 		default: edge_mask_reg_512p7[85] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100111,
11'b1111101000,
11'b10010000100,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10110010011,
11'b10110010100,
11'b10110100011,
11'b10110100100,
11'b10110110011,
11'b10110110100,
11'b10111000011,
11'b10111000100,
11'b10111010011,
11'b10111010100: edge_mask_reg_512p7[86] <= 1'b1;
 		default: edge_mask_reg_512p7[86] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111010110,
11'b111010111,
11'b111011000,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010111,
11'b10010000100,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000011,
11'b10011000100,
11'b10110010011,
11'b10110010100,
11'b10110100011,
11'b10110100100,
11'b10110110011,
11'b10110110100,
11'b10111000011,
11'b10111000100: edge_mask_reg_512p7[87] <= 1'b1;
 		default: edge_mask_reg_512p7[87] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[88] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111010110,
11'b111010111,
11'b111011000,
11'b1011010111,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111110111,
11'b10011110101,
11'b10011110110,
11'b10111110100,
11'b10111110101,
11'b10111110110,
11'b11011110100,
11'b11011110101,
11'b11111110101: edge_mask_reg_512p7[89] <= 1'b1;
 		default: edge_mask_reg_512p7[89] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100110,
11'b10010100111,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100110,
11'b10110100111,
11'b11001100110,
11'b11001100111,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11010000110,
11'b11010000111,
11'b11010010110,
11'b11010010111,
11'b11010100110,
11'b11010100111,
11'b11101100110,
11'b11101100111,
11'b11101110110,
11'b11101110111,
11'b11110000110,
11'b11110000111,
11'b11110010110,
11'b11110010111,
11'b11110100110,
11'b11110100111: edge_mask_reg_512p7[90] <= 1'b1;
 		default: edge_mask_reg_512p7[90] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010100,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101001,
11'b1011101010,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100100,
11'b1111101001,
11'b1111101010,
11'b10010110101,
11'b10010110110,
11'b10010111010,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011100100: edge_mask_reg_512p7[91] <= 1'b1;
 		default: edge_mask_reg_512p7[91] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011100110,
11'b10011100111,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111100110,
11'b10111100111,
11'b10111110110,
11'b10111110111,
11'b11011100110,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111110101,
11'b11111110110: edge_mask_reg_512p7[92] <= 1'b1;
 		default: edge_mask_reg_512p7[92] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111010110,
11'b10111010111,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111100101,
11'b11111100110,
11'b11111110101,
11'b11111110110: edge_mask_reg_512p7[93] <= 1'b1;
 		default: edge_mask_reg_512p7[93] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011101001: edge_mask_reg_512p7[94] <= 1'b1;
 		default: edge_mask_reg_512p7[94] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101001,
11'b1010101010,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000111,
11'b10110001000,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11010000111,
11'b11010001000,
11'b11101010110,
11'b11101100110,
11'b11101100111,
11'b11101110110,
11'b11101110111: edge_mask_reg_512p7[95] <= 1'b1;
 		default: edge_mask_reg_512p7[95] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111011,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010011001,
11'b10101100111,
11'b10101101000,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10101111010,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110001010,
11'b10110011000,
11'b10110011001,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11010000111,
11'b11010001000,
11'b11010001001,
11'b11010011000,
11'b11010011001,
11'b11101100110,
11'b11101100111,
11'b11101110110,
11'b11101110111,
11'b11101111000,
11'b11101111001,
11'b11110000111,
11'b11110001000,
11'b11110001001: edge_mask_reg_512p7[96] <= 1'b1;
 		default: edge_mask_reg_512p7[96] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001010,
11'b111001011,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001010,
11'b1011001011,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10101100111,
11'b10101101000,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100111,
11'b10110101000,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11010000110,
11'b11010000111,
11'b11010001000,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010100111,
11'b11101100110,
11'b11101100111,
11'b11101110110,
11'b11101110111,
11'b11110000110: edge_mask_reg_512p7[97] <= 1'b1;
 		default: edge_mask_reg_512p7[97] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b11010100110,
11'b11010100111,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000101,
11'b11011000110,
11'b11011000111,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11110110101,
11'b11110110110,
11'b11110110111,
11'b11111000101,
11'b11111000110,
11'b11111010101,
11'b11111010110: edge_mask_reg_512p7[98] <= 1'b1;
 		default: edge_mask_reg_512p7[98] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101010,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111101010,
11'b1111101011,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111001010,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11010111001,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011001001,
11'b11110101000,
11'b11110110110,
11'b11110110111,
11'b11110111000,
11'b11110111001,
11'b11111000110,
11'b11111000111,
11'b11111001000,
11'b11111001001: edge_mask_reg_512p7[99] <= 1'b1;
 		default: edge_mask_reg_512p7[99] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b11010100110,
11'b11010100111,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000101,
11'b11011000110,
11'b11011000111,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011100101,
11'b11011100110,
11'b11110110110,
11'b11110110111,
11'b11111000101,
11'b11111000110: edge_mask_reg_512p7[100] <= 1'b1;
 		default: edge_mask_reg_512p7[100] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000111,
11'b10011001000,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b11010100110,
11'b11010100111,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000101,
11'b11011000110,
11'b11011000111,
11'b11110110101,
11'b11110110110,
11'b11110110111,
11'b11111000110: edge_mask_reg_512p7[101] <= 1'b1;
 		default: edge_mask_reg_512p7[101] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011001,
11'b1111011010,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000111,
11'b10011001000,
11'b10101110111,
11'b10101111000,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000111,
11'b10111001000,
11'b11001110111,
11'b11001111000,
11'b11010000110,
11'b11010000111,
11'b11010001000,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000110,
11'b11011000111,
11'b11101110111,
11'b11101111000,
11'b11110000110,
11'b11110000111,
11'b11110001000,
11'b11110010110,
11'b11110010111,
11'b11110011000,
11'b11110100110,
11'b11110100111,
11'b11110101000,
11'b11110110110,
11'b11110110111,
11'b11111000110: edge_mask_reg_512p7[102] <= 1'b1;
 		default: edge_mask_reg_512p7[102] <= 1'b0;
 	endcase

    case({x,y,z})
11'b101011100,
11'b110011100,
11'b110101100,
11'b1000111100,
11'b1001001100,
11'b1001001101,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011100,
11'b1010011101,
11'b1010101100,
11'b1010101101,
11'b1010111100,
11'b1010111101,
11'b1101001100,
11'b1101001101,
11'b1101011100,
11'b1101011101,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101100,
11'b1110101101,
11'b1110111101,
11'b1111001101,
11'b10001101010,
11'b10001101011,
11'b10001101100,
11'b10001101101,
11'b10001101110,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10001111101,
11'b10001111110,
11'b10010001010,
11'b10010001011,
11'b10010001100,
11'b10010001101,
11'b10010001110,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10010011101,
11'b10010011110,
11'b10101101001,
11'b10101101010,
11'b10101101011,
11'b10101101100,
11'b10101111001,
11'b10101111010,
11'b10101111011,
11'b10101111100,
11'b10101111101,
11'b10110001001,
11'b10110001010,
11'b10110001011,
11'b10110001100,
11'b10110011010,
11'b10110011011,
11'b10110011100,
11'b11001101001,
11'b11001101010,
11'b11001101011,
11'b11001111001,
11'b11001111010,
11'b11001111011,
11'b11001111100,
11'b11010001001,
11'b11010001010,
11'b11010001011,
11'b11010001100,
11'b11010011010,
11'b11010011011,
11'b11010011100,
11'b11101111001,
11'b11101111010,
11'b11101111011,
11'b11110001001,
11'b11110001010,
11'b11110001011,
11'b11110011010,
11'b11110011011: edge_mask_reg_512p7[103] <= 1'b1;
 		default: edge_mask_reg_512p7[103] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000101001,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10000111010,
11'b10000111011,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10100010101,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000110,
11'b10101000111: edge_mask_reg_512p7[104] <= 1'b1;
 		default: edge_mask_reg_512p7[104] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000101: edge_mask_reg_512p7[105] <= 1'b1;
 		default: edge_mask_reg_512p7[105] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b101000110,
11'b101000111,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010011,
11'b1001010100,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100011,
11'b1110101000,
11'b10001010011,
11'b10001100011,
11'b10001110011,
11'b10001110100,
11'b10010000011,
11'b10010000100,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p7[106] <= 1'b1;
 		default: edge_mask_reg_512p7[106] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[107] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[108] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[109] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[110] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[111] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b10010010110,
11'b10010010111,
11'b10010100110,
11'b10010100111,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000111,
11'b10011001000,
11'b10011010111,
11'b10011011000,
11'b10110010110,
11'b10110010111,
11'b10110100110,
11'b10110100111,
11'b10110110110,
11'b10110110111,
11'b10111000111,
11'b10111001000,
11'b10111010111,
11'b10111011000,
11'b11010010110,
11'b11010010111,
11'b11010100110,
11'b11010100111,
11'b11010110111,
11'b11011000111,
11'b11011010111,
11'b11110010110,
11'b11110010111,
11'b11110100110,
11'b11110100111,
11'b11110110111,
11'b11111000111,
11'b11111010111: edge_mask_reg_512p7[112] <= 1'b1;
 		default: edge_mask_reg_512p7[112] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110111,
11'b10010111000,
11'b10011000111,
11'b10011001000,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110111,
11'b10110111000,
11'b10111000111,
11'b10111001000,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110111,
11'b11010111000,
11'b11011000111,
11'b11011001000,
11'b11110010110,
11'b11110010111,
11'b11110100110,
11'b11110100111,
11'b11110101000,
11'b11110110111,
11'b11110111000,
11'b11111000111,
11'b11111001000: edge_mask_reg_512p7[113] <= 1'b1;
 		default: edge_mask_reg_512p7[113] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000011000,
11'b1000011001: edge_mask_reg_512p7[114] <= 1'b1;
 		default: edge_mask_reg_512p7[114] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000011000,
11'b1000011001: edge_mask_reg_512p7[115] <= 1'b1;
 		default: edge_mask_reg_512p7[115] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111001,
11'b1000111010,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100111001,
11'b1100111010,
11'b10000010111,
11'b10000011000,
11'b10100000110,
11'b10100000111,
11'b10100001000,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b11000000101,
11'b11000000110,
11'b11000000111,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11100000101,
11'b11100000110,
11'b11100000111,
11'b11100010101,
11'b11100010110,
11'b11100010111: edge_mask_reg_512p7[116] <= 1'b1;
 		default: edge_mask_reg_512p7[116] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000011000,
11'b1000011001,
11'b1000101001,
11'b1100011000,
11'b1100011001,
11'b10100000110,
11'b10100000111,
11'b11000000110: edge_mask_reg_512p7[117] <= 1'b1;
 		default: edge_mask_reg_512p7[117] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001001,
11'b1101001010,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000110111,
11'b10100000110,
11'b10100000111,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b11000000101,
11'b11000000110,
11'b11000000111,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11000100101,
11'b11000100110,
11'b11000100111,
11'b11000110101,
11'b11000110110,
11'b11100000101: edge_mask_reg_512p7[118] <= 1'b1;
 		default: edge_mask_reg_512p7[118] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010101000,
11'b10010101001,
11'b10010111000,
11'b10010111001,
11'b10011001000,
11'b10011001001,
11'b10011011000,
11'b10011011001,
11'b10011101000,
11'b10011101001,
11'b10110101000,
11'b10110101001,
11'b10110111000,
11'b10110111001,
11'b10111001000,
11'b10111001001,
11'b10111011000,
11'b10111011001,
11'b10111101000,
11'b10111101001,
11'b11010101000,
11'b11010101001,
11'b11010111000,
11'b11010111001,
11'b11011001000,
11'b11011001001,
11'b11011011000,
11'b11011011001,
11'b11011101000,
11'b11011101001,
11'b11110100111,
11'b11110101000,
11'b11110110111,
11'b11110111000,
11'b11110111001,
11'b11111001000,
11'b11111001001,
11'b11111011000,
11'b11111011001,
11'b11111101000,
11'b11111101001: edge_mask_reg_512p7[119] <= 1'b1;
 		default: edge_mask_reg_512p7[119] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[120] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[121] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[122] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[123] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101011,
11'b100101010,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b1000011001,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011011,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10000011011,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000101011,
11'b10000111000,
11'b10000111001,
11'b10000111011,
11'b10100000110,
11'b10100000111,
11'b10100001000,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100011001,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100101001,
11'b10100110111,
11'b10100111000,
11'b10100111001,
11'b11000000110,
11'b11000001000,
11'b11000010110,
11'b11000010111,
11'b11000011000,
11'b11000100110,
11'b11000100111,
11'b11000101000,
11'b11000110111,
11'b11000111000: edge_mask_reg_512p7[124] <= 1'b1;
 		default: edge_mask_reg_512p7[124] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011011,
11'b100101001,
11'b100101010,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10000011011,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000101010,
11'b10000101011,
11'b10100000111,
11'b10100001000,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100110,
11'b10100100111: edge_mask_reg_512p7[125] <= 1'b1;
 		default: edge_mask_reg_512p7[125] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111010,
11'b11001010,
11'b110111011,
11'b110111100,
11'b111001010,
11'b111001011,
11'b111011010,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101010,
11'b1111001011,
11'b1111001100,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111111000,
11'b1111111001,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101011,
11'b10011111000,
11'b10011111001,
11'b10011111010,
11'b10111101000,
11'b10111101001,
11'b10111111000,
11'b10111111001,
11'b10111111010,
11'b11011101000,
11'b11011101001,
11'b11011111000,
11'b11011111001,
11'b11111100111,
11'b11111101000,
11'b11111110111,
11'b11111111000,
11'b11111111001: edge_mask_reg_512p7[126] <= 1'b1;
 		default: edge_mask_reg_512p7[126] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1100111010,
11'b1100111011,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010011001,
11'b10101010111,
11'b10101011000,
11'b10101011001,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10101111010,
11'b10110001000,
11'b10110001001,
11'b10110001010,
11'b10110011001,
11'b11001010111,
11'b11001011000,
11'b11001100111,
11'b11001101000,
11'b11001101001,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11010001000,
11'b11010001001,
11'b11010011000,
11'b11010011001,
11'b11101010111,
11'b11101011000,
11'b11101100111,
11'b11101101000,
11'b11101101001,
11'b11101110111,
11'b11101111000,
11'b11101111001,
11'b11110001000,
11'b11110001001: edge_mask_reg_512p7[127] <= 1'b1;
 		default: edge_mask_reg_512p7[127] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000111,
11'b11001000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10110100011,
11'b10110100100,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111010011,
11'b10111010100,
11'b11010110100,
11'b11011000100,
11'b11011010100: edge_mask_reg_512p7[128] <= 1'b1;
 		default: edge_mask_reg_512p7[128] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100111,
11'b1101101000,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10100010100,
11'b10100010101,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110100,
11'b10100110101,
11'b10101000100,
11'b10101000101,
11'b10101010100,
11'b10101010101,
11'b11000010100,
11'b11000010101,
11'b11000100100,
11'b11000100101,
11'b11000110100,
11'b11000110101,
11'b11001000100,
11'b11001000101: edge_mask_reg_512p7[129] <= 1'b1;
 		default: edge_mask_reg_512p7[129] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000111,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110100,
11'b10000110101,
11'b10100010100,
11'b10100010101,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b11000010100,
11'b11000010101,
11'b11000100100,
11'b11000110100: edge_mask_reg_512p7[130] <= 1'b1;
 		default: edge_mask_reg_512p7[130] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110111,
11'b1100111000,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10100010100,
11'b10100010101,
11'b10100100100,
11'b10100100101,
11'b11000000101,
11'b11000010100,
11'b11000010101,
11'b11100000101,
11'b11100010100: edge_mask_reg_512p7[131] <= 1'b1;
 		default: edge_mask_reg_512p7[131] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110111,
11'b1100111000,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10100010100,
11'b10100010101,
11'b10100100100,
11'b10100100101,
11'b11000010100,
11'b11000010101: edge_mask_reg_512p7[132] <= 1'b1;
 		default: edge_mask_reg_512p7[132] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110111,
11'b1100111000,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10100010100,
11'b10100010101,
11'b10100100100,
11'b10100100101,
11'b11000010100,
11'b11000010101,
11'b11100010100: edge_mask_reg_512p7[133] <= 1'b1;
 		default: edge_mask_reg_512p7[133] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110101000,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100111,
11'b10011101000,
11'b10110110110,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100111,
11'b10111101000,
11'b11011000110,
11'b11011000111,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100111,
11'b11011101000,
11'b11111000110,
11'b11111000111,
11'b11111010110,
11'b11111010111,
11'b11111011000,
11'b11111100111,
11'b11111101000: edge_mask_reg_512p7[134] <= 1'b1;
 		default: edge_mask_reg_512p7[134] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111010,
11'b1010111011,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111010,
11'b1110111011,
11'b10001111001,
11'b10001111010,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10101111000,
11'b10101111001,
11'b10101111010,
11'b10110001000,
11'b10110001001,
11'b10110001010,
11'b10110011000,
11'b10110011001,
11'b10110011010,
11'b11001111000,
11'b11001111001,
11'b11010001000,
11'b11010001001,
11'b11010011000,
11'b11010011001,
11'b11101111000,
11'b11101111001,
11'b11110001000,
11'b11110001001,
11'b11110011000,
11'b11110011001: edge_mask_reg_512p7[135] <= 1'b1;
 		default: edge_mask_reg_512p7[135] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[136] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[137] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[138] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[139] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[140] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[141] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011011,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001001,
11'b1101001010,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10100000110,
11'b10100000111,
11'b10100001000,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b11000000101,
11'b11000000110,
11'b11000000111,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11000100101,
11'b11000100110,
11'b11000100111: edge_mask_reg_512p7[142] <= 1'b1;
 		default: edge_mask_reg_512p7[142] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[143] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100111,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000110,
11'b10001000111,
11'b10100000111,
11'b10100001000,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b11000000111,
11'b11000010110,
11'b11000010111,
11'b11000011000,
11'b11000100101,
11'b11000100110,
11'b11000100111,
11'b11000101000,
11'b11000110101,
11'b11000110110,
11'b11000110111,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010101,
11'b11001010110,
11'b11100000111,
11'b11100010110,
11'b11100010111,
11'b11100011000,
11'b11100100101,
11'b11100100110,
11'b11100100111,
11'b11100101000,
11'b11100110101,
11'b11100110110,
11'b11100110111,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101010110: edge_mask_reg_512p7[144] <= 1'b1;
 		default: edge_mask_reg_512p7[144] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101010,
11'b10101011,
11'b10111011,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111011,
11'b101111100,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b1000101011,
11'b1000111011,
11'b1000111100,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1100101100,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b10001001000,
11'b10001001001,
11'b10001001100,
11'b10001001101,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001011010,
11'b10001011100,
11'b10001011101,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101100,
11'b10001101101,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001011,
11'b10010001100,
11'b10101010111,
11'b10101011000,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000111,
11'b10110001000,
11'b11001010111,
11'b11001100111,
11'b11001101000,
11'b11001110111,
11'b11001111000,
11'b11010000111,
11'b11010001000: edge_mask_reg_512p7[145] <= 1'b1;
 		default: edge_mask_reg_512p7[145] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101010,
11'b10101011,
11'b10111010,
11'b10111011,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001010,
11'b111001011,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001011,
11'b1011001100,
11'b1011011011,
11'b1011011100,
11'b1101001011,
11'b1101001100,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001011,
11'b1111001100,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010001100,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010101100,
11'b10101101000,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110011010,
11'b10110101000,
11'b10110101001,
11'b11001110111,
11'b11001111000,
11'b11010000111,
11'b11010001000,
11'b11010001001,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11110000111,
11'b11110001000,
11'b11110010111,
11'b11110011000,
11'b11110100111,
11'b11110101000: edge_mask_reg_512p7[146] <= 1'b1;
 		default: edge_mask_reg_512p7[146] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101010,
11'b10101011,
11'b10111011,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b1000101011,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1100101011,
11'b1100101100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001011011,
11'b10001011100,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001101100,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001011,
11'b10010001100,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000111,
11'b10110001000,
11'b11001000110,
11'b11001010110,
11'b11001010111,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11010000111,
11'b11010001000: edge_mask_reg_512p7[147] <= 1'b1;
 		default: edge_mask_reg_512p7[147] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101001,
11'b10101010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000010111,
11'b1000011000,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110011000,
11'b10000100101,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10100100101,
11'b10100100110,
11'b10100110101,
11'b10100110110,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100110,
11'b10101100111,
11'b10101110110,
11'b10101110111,
11'b11000100101,
11'b11000110101,
11'b11000110110,
11'b11001000101,
11'b11001000110,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110110,
11'b11001110111,
11'b11100110101,
11'b11100110110,
11'b11101000101,
11'b11101000110,
11'b11101010101,
11'b11101010110,
11'b11101010111,
11'b11101100110,
11'b11101100111,
11'b11101110110,
11'b11101110111: edge_mask_reg_512p7[148] <= 1'b1;
 		default: edge_mask_reg_512p7[148] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101001,
11'b10101010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110011000,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10100110110,
11'b10100110111,
11'b10101000110,
11'b10101000111,
11'b10101010110,
11'b10101010111,
11'b10101100110,
11'b10101100111,
11'b10101110110,
11'b10101110111,
11'b11000110110,
11'b11000110111,
11'b11001000110,
11'b11001000111,
11'b11001010110,
11'b11001010111,
11'b11001100110,
11'b11001100111,
11'b11001110110,
11'b11001110111,
11'b11100110110,
11'b11100110111,
11'b11101000110,
11'b11101000111,
11'b11101010110,
11'b11101010111,
11'b11101100110,
11'b11101100111,
11'b11101110110,
11'b11101110111: edge_mask_reg_512p7[149] <= 1'b1;
 		default: edge_mask_reg_512p7[149] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101001,
11'b10101010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1100110111,
11'b1100111000,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110011000,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010110,
11'b10001010111,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10100110110,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100110,
11'b10101100111,
11'b10101110110,
11'b10101110111,
11'b11001000101,
11'b11001000110,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001110110,
11'b11001110111,
11'b11101000101,
11'b11101000110,
11'b11101010101,
11'b11101010110,
11'b11101010111,
11'b11101100110,
11'b11101100111,
11'b11101110110,
11'b11101110111: edge_mask_reg_512p7[150] <= 1'b1;
 		default: edge_mask_reg_512p7[150] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101001,
11'b10101010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000010111,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110011000,
11'b10000110110,
11'b10000110111,
11'b10001000110,
11'b10001000111,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10100110110,
11'b10100110111,
11'b10101000110,
11'b10101000111,
11'b10101010110,
11'b10101010111,
11'b10101100110,
11'b10101100111,
11'b10101110110,
11'b10101110111,
11'b11000110101,
11'b11000110110,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010110,
11'b11001010111,
11'b11001100110,
11'b11001100111,
11'b11001110110,
11'b11001110111,
11'b11100110101,
11'b11100110110,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101010110,
11'b11101010111,
11'b11101100110,
11'b11101100111,
11'b11101110110,
11'b11101110111: edge_mask_reg_512p7[151] <= 1'b1;
 		default: edge_mask_reg_512p7[151] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000110,
11'b10010000111,
11'b10010010110,
11'b10010010111,
11'b10101100110,
11'b10101100111,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b11001100110,
11'b11001100111,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010101,
11'b11010010110,
11'b11101100110,
11'b11101100111,
11'b11101110110,
11'b11101110111,
11'b11110000101,
11'b11110000110,
11'b11110000111,
11'b11110010101,
11'b11110010110: edge_mask_reg_512p7[152] <= 1'b1;
 		default: edge_mask_reg_512p7[152] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101001,
11'b10101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10101010111,
11'b10101011000,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b11001010111,
11'b11001011000,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11101010111,
11'b11101011000,
11'b11101100110,
11'b11101100111,
11'b11101101000,
11'b11101110110,
11'b11101110111,
11'b11101111000: edge_mask_reg_512p7[153] <= 1'b1;
 		default: edge_mask_reg_512p7[153] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b10001011001,
11'b10001011010,
11'b10001011011,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10101011001,
11'b10101011010,
11'b10101101000,
11'b10101101001,
11'b10101101010,
11'b10101101011,
11'b10101111001,
11'b10101111010,
11'b10101111011,
11'b11001011000,
11'b11001011001,
11'b11001011010,
11'b11001101000,
11'b11001101001,
11'b11001101010,
11'b11001101011,
11'b11001111001,
11'b11001111010,
11'b11001111011,
11'b11101011000,
11'b11101011001,
11'b11101011010,
11'b11101101000,
11'b11101101001,
11'b11101101010,
11'b11101101011,
11'b11101111001,
11'b11101111010,
11'b11101111011: edge_mask_reg_512p7[154] <= 1'b1;
 		default: edge_mask_reg_512p7[154] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[155] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[156] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10011010101,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10011110111,
11'b10011111000,
11'b10011111001,
11'b10111000101,
11'b10111000110,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b10111111001,
11'b11011000101,
11'b11011000110,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011101000,
11'b11011110110,
11'b11011110111,
11'b11011111000,
11'b11111000101,
11'b11111000110,
11'b11111010101,
11'b11111010110,
11'b11111010111,
11'b11111100110,
11'b11111100111,
11'b11111101000,
11'b11111110110,
11'b11111110111,
11'b11111111000: edge_mask_reg_512p7[157] <= 1'b1;
 		default: edge_mask_reg_512p7[157] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100100111,
11'b100101000,
11'b100101001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b10000010111,
11'b10000011000,
11'b10100000111,
11'b10100001000,
11'b10100001001,
11'b10100010111,
11'b10100011000,
11'b11000000111,
11'b11000001000,
11'b11000001001,
11'b11000010111,
11'b11000011000,
11'b11100000111,
11'b11100001000,
11'b11100001001,
11'b11100010111,
11'b11100011000: edge_mask_reg_512p7[158] <= 1'b1;
 		default: edge_mask_reg_512p7[158] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100111000,
11'b1100111001,
11'b10000011000,
11'b10000011001,
11'b10100001000,
11'b10100001001,
11'b10100011000,
11'b10100011001,
11'b11000001000,
11'b11000001001,
11'b11000011000,
11'b11000011001,
11'b11100000111,
11'b11100001000,
11'b11100001001,
11'b11100011000,
11'b11100011001: edge_mask_reg_512p7[159] <= 1'b1;
 		default: edge_mask_reg_512p7[159] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1100100111,
11'b1100101000,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110111,
11'b1101111000,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10100110100,
11'b10100110101,
11'b10101000100,
11'b10101000101,
11'b10101010100,
11'b10101010101,
11'b10101100100,
11'b10101100101,
11'b11000110100,
11'b11000110101,
11'b11001000100,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11001100101,
11'b11101000100,
11'b11101010100: edge_mask_reg_512p7[160] <= 1'b1;
 		default: edge_mask_reg_512p7[160] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110111,
11'b1101111000,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b11000010101,
11'b11000100100,
11'b11000100101,
11'b11000110100,
11'b11000110101,
11'b11001000100,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11001100101,
11'b11100100100,
11'b11100110100,
11'b11101000100,
11'b11101010100: edge_mask_reg_512p7[161] <= 1'b1;
 		default: edge_mask_reg_512p7[161] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110111,
11'b1101111000,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10100010100,
11'b10100010101,
11'b10100100100,
11'b10100100101,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10101000100,
11'b10101000101,
11'b10101010100,
11'b10101010101,
11'b10101100100,
11'b10101100101,
11'b11000010100,
11'b11000010101,
11'b11000100100,
11'b11000100101,
11'b11000110100,
11'b11000110101,
11'b11001000100,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11001100101,
11'b11100100100,
11'b11100110100,
11'b11101000100,
11'b11101010100: edge_mask_reg_512p7[162] <= 1'b1;
 		default: edge_mask_reg_512p7[162] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[163] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101011,
11'b10111011,
11'b101001011,
11'b101001100,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b101111011,
11'b101111100,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b111001011,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001011,
11'b1011001100,
11'b1011011011,
11'b1011011100,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b1111011011,
11'b1111011100,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001101100,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10001111101,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010001100,
11'b10010001101,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10010011101,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010101011,
11'b10010101100,
11'b10010111000,
11'b10010111001,
11'b10101101000,
11'b10101101001,
11'b10101101010,
11'b10101111000,
11'b10101111001,
11'b10101111010,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110001010,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110011010,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110111000,
11'b11001111000,
11'b11001111001,
11'b11010000111,
11'b11010001000,
11'b11010001001,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010100111,
11'b11010101000,
11'b11101111000,
11'b11101111001,
11'b11110001000,
11'b11110001001,
11'b11110011000: edge_mask_reg_512p7[164] <= 1'b1;
 		default: edge_mask_reg_512p7[164] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[165] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[166] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[167] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[168] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[169] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[170] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101001,
11'b10101010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010011000,
11'b1010011001,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110011000,
11'b1110011001,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010111,
11'b10001011000,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100111,
11'b11001101000,
11'b11001101001,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11100110110,
11'b11100110111,
11'b11101000110,
11'b11101000111,
11'b11101001000,
11'b11101010110,
11'b11101010111,
11'b11101011000,
11'b11101100111,
11'b11101101000,
11'b11101110111,
11'b11101111000,
11'b11110000111,
11'b11110001000: edge_mask_reg_512p7[171] <= 1'b1;
 		default: edge_mask_reg_512p7[171] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011100110,
11'b1011100111,
11'b1111100110,
11'b11011110101,
11'b11111110101: edge_mask_reg_512p7[172] <= 1'b1;
 		default: edge_mask_reg_512p7[172] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011100110,
11'b1011100111,
11'b1111100110,
11'b11011110101,
11'b11111110101: edge_mask_reg_512p7[173] <= 1'b1;
 		default: edge_mask_reg_512p7[173] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110011000,
11'b1110011001,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111111000,
11'b1111111001,
11'b10010100100,
11'b10010100101,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011010111,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10110100100,
11'b10110100101,
11'b10110110011,
11'b10110110100,
11'b10110110101,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111000110,
11'b10111010011,
11'b10111010100,
11'b10111010101,
11'b10111010110,
11'b10111100011,
11'b10111100100,
11'b10111100101,
11'b10111100110,
11'b10111110100,
11'b10111110101: edge_mask_reg_512p7[174] <= 1'b1;
 		default: edge_mask_reg_512p7[174] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101010,
11'b1111011011,
11'b1111011100,
11'b1111101010,
11'b1111101011,
11'b1111111000,
11'b1111111001,
11'b10011111000,
11'b10011111001,
11'b10111110111,
11'b10111111000,
11'b10111111001,
11'b11011111000,
11'b11011111001: edge_mask_reg_512p7[175] <= 1'b1;
 		default: edge_mask_reg_512p7[175] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001010,
11'b1110001011,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001011010,
11'b10001011011,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001110110,
11'b10001110111,
11'b10100110110,
11'b10100110111,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110111: edge_mask_reg_512p7[176] <= 1'b1;
 		default: edge_mask_reg_512p7[176] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011100,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101110101,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001001011,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011011,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101011,
11'b10100110110,
11'b10101000110,
11'b10101000111,
11'b10101010110,
11'b10101010111,
11'b10101100110,
11'b10101100111: edge_mask_reg_512p7[177] <= 1'b1;
 		default: edge_mask_reg_512p7[177] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[178] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[179] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[180] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[181] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[182] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[183] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b101111011,
11'b101111100,
11'b110001100,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111100,
11'b1101111101,
11'b10000100111,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10000111010,
11'b10000111100,
11'b10000111101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001001100,
11'b10001001101,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10100100111,
11'b10100101000,
11'b10100101001,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10100111001,
11'b10101000110,
11'b10101000111,
11'b10101001000: edge_mask_reg_512p7[184] <= 1'b1;
 		default: edge_mask_reg_512p7[184] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101011,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101100,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b10000100111,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10000111010,
11'b10000111100,
11'b10000111101,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001001010,
11'b10001001100,
11'b10001001101,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001011010,
11'b10001011100,
11'b10001011101,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101100,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111100,
11'b10100100111,
11'b10100101000,
11'b10100101001,
11'b10100110111,
11'b10100111000,
11'b10100111001,
11'b10101000111,
11'b10101001000,
11'b10101001001,
11'b10101010111,
11'b10101011000,
11'b10101011001,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101111000,
11'b10101111001,
11'b11000110111,
11'b11001000111,
11'b11001001000,
11'b11001010111,
11'b11001011000,
11'b11001011001,
11'b11001100111,
11'b11001101000,
11'b11001101001,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11101010111,
11'b11101100111,
11'b11101101000: edge_mask_reg_512p7[185] <= 1'b1;
 		default: edge_mask_reg_512p7[185] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[186] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010111,
11'b1001011000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b10100110100,
11'b10100110101,
11'b11000000101,
11'b11000000110,
11'b11000010100,
11'b11000010101,
11'b11000100100,
11'b11000100101,
11'b11000110100,
11'b11000110101,
11'b11100000101,
11'b11100010100,
11'b11100100100: edge_mask_reg_512p7[187] <= 1'b1;
 		default: edge_mask_reg_512p7[187] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100101000,
11'b100101001,
11'b100101010,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100101000,
11'b1100101001,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10100010101,
11'b10100010110,
11'b11000000101,
11'b11000000110,
11'b11000010101,
11'b11100000101: edge_mask_reg_512p7[188] <= 1'b1;
 		default: edge_mask_reg_512p7[188] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10001010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1100011000,
11'b1100011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101101000,
11'b1101101001,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100101,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101100101,
11'b11000100100,
11'b11000100101,
11'b11000100110,
11'b11000110100,
11'b11000110101,
11'b11000110110,
11'b11001000100,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11100100100,
11'b11100100101,
11'b11100110100,
11'b11100110101,
11'b11101000100,
11'b11101000101,
11'b11101010100: edge_mask_reg_512p7[189] <= 1'b1;
 		default: edge_mask_reg_512p7[189] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b10000110101,
11'b10000110110,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10100110101,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000100,
11'b10110000101,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11010000101,
11'b11101000100,
11'b11101000101,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101,
11'b11101110100: edge_mask_reg_512p7[190] <= 1'b1;
 		default: edge_mask_reg_512p7[190] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111001,
11'b1000111010,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100111001,
11'b1100111010,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10100000110,
11'b10100000111,
11'b10100001000,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b11000000101,
11'b11000000110,
11'b11000000111,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11100000101,
11'b11100000110,
11'b11100000111,
11'b11100010101,
11'b11100010110,
11'b11100010111: edge_mask_reg_512p7[191] <= 1'b1;
 		default: edge_mask_reg_512p7[191] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[192] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[193] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[194] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100101010,
11'b1000011001,
11'b1000101001,
11'b1000101010,
11'b1100011001,
11'b1100011010,
11'b1100101001,
11'b1100101010,
11'b10000011000,
11'b10100000111,
11'b10100001000,
11'b10100011000,
11'b11000000110,
11'b11000000111,
11'b11000001000,
11'b11000010110,
11'b11000010111,
11'b11100000110,
11'b11100000111,
11'b11100001000,
11'b11100010110,
11'b11100010111: edge_mask_reg_512p7[195] <= 1'b1;
 		default: edge_mask_reg_512p7[195] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[196] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011011,
11'b1101010,
11'b1101011,
11'b100111011,
11'b101001011,
11'b101001100,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b101111100,
11'b1000101011,
11'b1000111011,
11'b1000111100,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1100011010,
11'b1100011011,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b10000011010,
11'b10000011011,
11'b10000101010,
11'b10000101011,
11'b10000101100,
11'b10000111010,
11'b10000111011,
11'b10000111100,
11'b10000111101,
11'b10001001010,
11'b10001001011,
11'b10100011010,
11'b10100011011,
11'b10100101001,
11'b10100101010,
11'b10100101011,
11'b10100111001,
11'b10100111010,
11'b10100111011,
11'b10101001001,
11'b10101001010,
11'b10101001011,
11'b11000001010,
11'b11000001011,
11'b11000011001,
11'b11000011010,
11'b11000011011,
11'b11000101001,
11'b11000101010,
11'b11000101011,
11'b11000111001,
11'b11000111010,
11'b11000111011,
11'b11001001001,
11'b11001001010,
11'b11100001001,
11'b11100001010,
11'b11100001011,
11'b11100011001,
11'b11100011010,
11'b11100011011,
11'b11100101001,
11'b11100101010,
11'b11100101011,
11'b11100111001,
11'b11100111010,
11'b11101001010: edge_mask_reg_512p7[197] <= 1'b1;
 		default: edge_mask_reg_512p7[197] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001010,
11'b1011010,
11'b1011011,
11'b1101011,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101100,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000101,
11'b1001000110,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011011,
11'b1001011100,
11'b1100011010,
11'b1100011011,
11'b1100100100,
11'b1100100101,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100110100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011011,
11'b1101011100,
11'b10000011011,
11'b10000101011,
11'b10000101100,
11'b10000111100: edge_mask_reg_512p7[198] <= 1'b1;
 		default: edge_mask_reg_512p7[198] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001011,
11'b10011011,
11'b10101011,
11'b10111011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b111001011,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101010,
11'b1110011100,
11'b1110011101,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10010111001,
11'b10010111010,
11'b10010111011,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011001100,
11'b10011001101,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011011100,
11'b10011011101,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101011,
11'b10011111000,
11'b10011111001,
11'b10011111010,
11'b10110111001,
11'b10110111010,
11'b10111001001,
11'b10111001010,
11'b10111011001,
11'b10111011010,
11'b10111101000,
11'b10111101001,
11'b10111101010,
11'b10111111000,
11'b10111111001,
11'b10111111010,
11'b11010111001,
11'b11011001001,
11'b11011001010,
11'b11011011001,
11'b11011011010,
11'b11011101001,
11'b11011101010,
11'b11011111001,
11'b11111001001,
11'b11111001010,
11'b11111011001,
11'b11111011010,
11'b11111101001,
11'b11111111001: edge_mask_reg_512p7[199] <= 1'b1;
 		default: edge_mask_reg_512p7[199] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[200] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[201] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[202] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1100111011,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b10001011000,
11'b10001011001,
11'b10001011010,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10101010111,
11'b10101011000,
11'b10101011001,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110001000,
11'b10110001001,
11'b10110011000,
11'b10110011001,
11'b11001010111,
11'b11001011000,
11'b11001100111,
11'b11001101000,
11'b11001101001,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11010001000,
11'b11010001001,
11'b11010011000,
11'b11010011001,
11'b11101011000,
11'b11101011001,
11'b11101101000,
11'b11101101001,
11'b11101111000,
11'b11101111001,
11'b11110001000,
11'b11110001001: edge_mask_reg_512p7[203] <= 1'b1;
 		default: edge_mask_reg_512p7[203] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111011,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1100111011,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101010,
11'b1110101011,
11'b10001011000,
11'b10001011001,
11'b10001011010,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10101010111,
11'b10101011000,
11'b10101011001,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110001000,
11'b10110001001,
11'b11001010111,
11'b11001011000,
11'b11001100111,
11'b11001101000,
11'b11001101001,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11010001000,
11'b11010001001,
11'b11101011000,
11'b11101011001,
11'b11101101000,
11'b11101101001,
11'b11101111000,
11'b11101111001,
11'b11110001000,
11'b11110001001: edge_mask_reg_512p7[204] <= 1'b1;
 		default: edge_mask_reg_512p7[204] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b1000010111,
11'b1000011000,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b10000010100,
11'b10000010101,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10100010100,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010100,
11'b10101010101,
11'b11000100100,
11'b11000110100,
11'b11001000100,
11'b11001000101,
11'b11001010100,
11'b11100110100,
11'b11101000100: edge_mask_reg_512p7[205] <= 1'b1;
 		default: edge_mask_reg_512p7[205] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000010111,
11'b1000011000,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10000010100,
11'b10000010101,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10100010100,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b11000100100,
11'b11000110100,
11'b11000110101,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11100100100,
11'b11100110100,
11'b11100110101,
11'b11101000100,
11'b11101000101,
11'b11101010101: edge_mask_reg_512p7[206] <= 1'b1;
 		default: edge_mask_reg_512p7[206] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011010,
11'b10011011,
11'b10101010,
11'b10101011,
11'b10111010,
11'b10111011,
11'b11001010,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001010,
11'b111001011,
11'b111011010,
11'b1010011100,
11'b1010011101,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101010,
11'b1110011100,
11'b1110011101,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111111001,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011001100,
11'b10011001101,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011011100,
11'b10011011101,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101011,
11'b10011101100,
11'b10011111000,
11'b10011111001,
11'b10011111010,
11'b10111001001,
11'b10111001010,
11'b10111001011,
11'b10111011000,
11'b10111011001,
11'b10111011010,
11'b10111011011,
11'b10111101000,
11'b10111101001,
11'b10111101010,
11'b10111101011,
11'b10111111000,
11'b10111111001,
11'b10111111010,
11'b11011001001,
11'b11011001010,
11'b11011011000,
11'b11011011001,
11'b11011011010,
11'b11011101000,
11'b11011101001,
11'b11011101010,
11'b11011111000,
11'b11011111001,
11'b11111001001,
11'b11111001010,
11'b11111011000,
11'b11111011001,
11'b11111011010,
11'b11111100111,
11'b11111101000,
11'b11111101001,
11'b11111101010,
11'b11111110111,
11'b11111111000,
11'b11111111001: edge_mask_reg_512p7[207] <= 1'b1;
 		default: edge_mask_reg_512p7[207] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111010,
11'b11001000,
11'b11001001,
11'b11001010,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111010100,
11'b1111010101,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111111000,
11'b1111111001,
11'b10011100100,
11'b10011100101: edge_mask_reg_512p7[208] <= 1'b1;
 		default: edge_mask_reg_512p7[208] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111010,
11'b10111011,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001011,
11'b1001001100,
11'b1001001101,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001011,
11'b1011001100,
11'b1101011100,
11'b1101011101,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101110101,
11'b1101110110,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110100100,
11'b1110100101,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b10001111101,
11'b10010001011,
11'b10010001100,
11'b10010001101,
11'b10010011011,
11'b10010011100,
11'b10010011101,
11'b10010101100,
11'b10010101101: edge_mask_reg_512p7[209] <= 1'b1;
 		default: edge_mask_reg_512p7[209] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[210] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[211] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[212] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[213] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[214] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[215] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101100101,
11'b101100110,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1101110110,
11'b1101110111,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100101,
11'b10010100110,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10011010101,
11'b10011010110,
11'b10011010111,
11'b10110000100,
11'b10110000101,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110101,
11'b10110110110,
11'b10111000101,
11'b10111000110,
11'b10111010101,
11'b10111010110,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11011000100,
11'b11011000101,
11'b11011000110,
11'b11011010100,
11'b11011010101,
11'b11011010110,
11'b11110000100,
11'b11110000101,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101,
11'b11110110100,
11'b11110110101,
11'b11110110110,
11'b11111000100,
11'b11111000101,
11'b11111000110,
11'b11111010100,
11'b11111010101,
11'b11111010110: edge_mask_reg_512p7[216] <= 1'b1;
 		default: edge_mask_reg_512p7[216] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101010110,
11'b101010111,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b111000101,
11'b111000110,
11'b111000111,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1011000110,
11'b1011000111,
11'b1101100110,
11'b1101100111,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110110110,
11'b1110110111,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100101,
11'b10010100110,
11'b10101110100,
11'b10101110101,
11'b10110000100,
11'b10110000101,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11101110100,
11'b11101110101,
11'b11110000100,
11'b11110000101,
11'b11110010100,
11'b11110010101,
11'b11110100100,
11'b11110100101: edge_mask_reg_512p7[217] <= 1'b1;
 		default: edge_mask_reg_512p7[217] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001101010,
11'b1001101011,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101001,
11'b1011101010,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111101001,
11'b1111101010,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010111000,
11'b10010111001,
11'b10011001000,
11'b10011001001,
11'b10110001000,
11'b10110001001,
11'b10110011000,
11'b10110011001,
11'b10110101000,
11'b10110101001,
11'b10110111000,
11'b10110111001,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b11010001000,
11'b11010001001,
11'b11010011000,
11'b11010011001,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11010110111,
11'b11010111000,
11'b11010111001,
11'b11011000111,
11'b11011001000,
11'b11110001000,
11'b11110001001,
11'b11110011000,
11'b11110011001,
11'b11110100111,
11'b11110101000,
11'b11110110111,
11'b11110111000,
11'b11111000111,
11'b11111001000: edge_mask_reg_512p7[218] <= 1'b1;
 		default: edge_mask_reg_512p7[218] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001010,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001010,
11'b111001011,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b10001100111,
11'b10001101000,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010101000,
11'b10010101001,
11'b10101100111,
11'b10101101000,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110101000,
11'b10110101001,
11'b11001100111,
11'b11001101000,
11'b11001110111,
11'b11001111000,
11'b11010000111,
11'b11010001000,
11'b11010001001,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010101000,
11'b11010101001,
11'b11101110110,
11'b11101110111,
11'b11101111000,
11'b11110000110,
11'b11110000111,
11'b11110001000,
11'b11110001001,
11'b11110010111,
11'b11110011000,
11'b11110011001,
11'b11110101000: edge_mask_reg_512p7[219] <= 1'b1;
 		default: edge_mask_reg_512p7[219] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001010,
11'b100111010,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001010,
11'b111001011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b10001010111,
11'b10001011000,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010101000,
11'b10010101001,
11'b10101010111,
11'b10101011000,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110101000,
11'b10110101001,
11'b11001010111,
11'b11001100111,
11'b11001101000,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11010000111,
11'b11010001000,
11'b11010001001,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010101000,
11'b11010101001,
11'b11101100111,
11'b11101101000,
11'b11101110111,
11'b11101111000,
11'b11110000111,
11'b11110001000,
11'b11110001001,
11'b11110010111,
11'b11110011000,
11'b11110011001,
11'b11110101000: edge_mask_reg_512p7[220] <= 1'b1;
 		default: edge_mask_reg_512p7[220] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000010111: edge_mask_reg_512p7[221] <= 1'b1;
 		default: edge_mask_reg_512p7[221] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111001000,
11'b1111001001,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011010100,
11'b10011010101,
11'b10011100100,
11'b10011100101: edge_mask_reg_512p7[222] <= 1'b1;
 		default: edge_mask_reg_512p7[222] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001001,
11'b1110001010,
11'b10001001001,
11'b10001001010,
11'b10001001011,
11'b10001011001,
11'b10001011010,
11'b10001011011,
11'b10001101001,
11'b10001101010,
11'b10101001001,
11'b10101001010,
11'b10101001011,
11'b10101011001,
11'b10101011010,
11'b10101011011,
11'b10101101001,
11'b10101101010,
11'b11001001001,
11'b11001001010,
11'b11001001011,
11'b11001011001,
11'b11001011010,
11'b11001011011,
11'b11001101001,
11'b11001101010,
11'b11101001001,
11'b11101001010,
11'b11101001011,
11'b11101011001,
11'b11101011010,
11'b11101011011,
11'b11101101000,
11'b11101101001,
11'b11101101010: edge_mask_reg_512p7[223] <= 1'b1;
 		default: edge_mask_reg_512p7[223] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001010,
11'b110001011,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b10001001010,
11'b10001001011,
11'b10001011010,
11'b10001011011,
11'b10001101010,
11'b10001101011,
11'b10101001010,
11'b10101001011,
11'b10101011010,
11'b10101011011,
11'b10101101010,
11'b10101101011,
11'b11001001010,
11'b11001001011,
11'b11001011010,
11'b11001011011,
11'b11001011100,
11'b11001101010,
11'b11001101011,
11'b11001101100,
11'b11101001010,
11'b11101001011,
11'b11101011001,
11'b11101011010,
11'b11101011011,
11'b11101011100,
11'b11101101010,
11'b11101101011,
11'b11101101100: edge_mask_reg_512p7[224] <= 1'b1;
 		default: edge_mask_reg_512p7[224] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[225] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111011,
11'b1110111100,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011011011,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101011,
11'b10011110101,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10011111001,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b10111111000: edge_mask_reg_512p7[226] <= 1'b1;
 		default: edge_mask_reg_512p7[226] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011101010,
11'b1111101001,
11'b1111101010,
11'b1111101011: edge_mask_reg_512p7[227] <= 1'b1;
 		default: edge_mask_reg_512p7[227] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011010,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110101,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111000110,
11'b10111000111,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111010101,
11'b11111010110,
11'b11111100101,
11'b11111100110: edge_mask_reg_512p7[228] <= 1'b1;
 		default: edge_mask_reg_512p7[228] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010101011,
11'b1010101100,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b10011000110,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011010111,
11'b10011011011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10011101010,
11'b10011101011,
11'b10011110101,
11'b10011110110,
11'b10011110111: edge_mask_reg_512p7[229] <= 1'b1;
 		default: edge_mask_reg_512p7[229] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011101010,
11'b1111101001,
11'b1111101010,
11'b1111101011: edge_mask_reg_512p7[230] <= 1'b1;
 		default: edge_mask_reg_512p7[230] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011101010,
11'b1111101001,
11'b1111101010,
11'b1111101011: edge_mask_reg_512p7[231] <= 1'b1;
 		default: edge_mask_reg_512p7[231] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011101010,
11'b1111101001,
11'b1111101010,
11'b1111101011: edge_mask_reg_512p7[232] <= 1'b1;
 		default: edge_mask_reg_512p7[232] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[233] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000111,
11'b1010001000,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b10000110100,
11'b10000110101,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10100110100,
11'b10100110101,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b11000110100,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101,
11'b11101000100,
11'b11101000101,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101: edge_mask_reg_512p7[234] <= 1'b1;
 		default: edge_mask_reg_512p7[234] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110110,
11'b1001110111,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10100000110,
11'b10100010101,
11'b10100010110,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100100,
11'b11000000101,
11'b11000000110,
11'b11000010101,
11'b11000010110,
11'b11000100100,
11'b11000100101,
11'b11000100110,
11'b11000110100,
11'b11000110101,
11'b11001000100,
11'b11001000101,
11'b11001010100,
11'b11100010100,
11'b11100010101,
11'b11100100100,
11'b11100100101,
11'b11100110100,
11'b11100110101,
11'b11101000100,
11'b11101010100: edge_mask_reg_512p7[235] <= 1'b1;
 		default: edge_mask_reg_512p7[235] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10000110100,
11'b10000110101,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10100110100,
11'b10100110101,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b11000110100,
11'b11001000100,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11101000100,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101,
11'b11101110100,
11'b11101110101,
11'b11110000101: edge_mask_reg_512p7[236] <= 1'b1;
 		default: edge_mask_reg_512p7[236] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110110,
11'b101110111,
11'b101111000,
11'b1000010111,
11'b1000011000,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110110,
11'b1001110111,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100100,
11'b11000100100,
11'b11000100101,
11'b11000110100,
11'b11000110101,
11'b11001000100,
11'b11001000101,
11'b11001010100,
11'b11100100100,
11'b11100100101,
11'b11100110100,
11'b11100110101,
11'b11101000100,
11'b11101000101,
11'b11101010100: edge_mask_reg_512p7[237] <= 1'b1;
 		default: edge_mask_reg_512p7[237] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b10000110100,
11'b10000110101,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10100110100,
11'b10100110101,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b11000110100,
11'b11001000100,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11001100101,
11'b11001110100,
11'b11001110101,
11'b11010000100: edge_mask_reg_512p7[238] <= 1'b1;
 		default: edge_mask_reg_512p7[238] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111011000,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10111000101,
11'b10111000110,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11011000101,
11'b11110000100,
11'b11110000101,
11'b11110000110,
11'b11110010100,
11'b11110010101,
11'b11110010110,
11'b11110100100,
11'b11110100101,
11'b11110100110,
11'b11110110100,
11'b11110110101,
11'b11110110110: edge_mask_reg_512p7[239] <= 1'b1;
 		default: edge_mask_reg_512p7[239] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111010,
11'b10111011,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001011,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001011,
11'b1011001100,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010001100,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10101010101,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110101000,
11'b11001110110,
11'b11001110111,
11'b11010000110,
11'b11010000111,
11'b11010010111: edge_mask_reg_512p7[240] <= 1'b1;
 		default: edge_mask_reg_512p7[240] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011011000,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b11010010101,
11'b11010010110,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11110010101,
11'b11110100100,
11'b11110100101,
11'b11110100110,
11'b11110110100,
11'b11110110101,
11'b11110110110: edge_mask_reg_512p7[241] <= 1'b1;
 		default: edge_mask_reg_512p7[241] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101010,
11'b10101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b1000101000,
11'b1000101011,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010010110,
11'b1010010111,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1100101011,
11'b1100101100,
11'b1100110111,
11'b1100111000,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101011,
11'b1110101100,
11'b10001001100,
11'b10001011011,
11'b10001011100,
11'b10001100101,
11'b10001101011,
11'b10001101100,
11'b10001110101,
11'b10001111011,
11'b10010001011: edge_mask_reg_512p7[242] <= 1'b1;
 		default: edge_mask_reg_512p7[242] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[243] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101001010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000100111,
11'b10000101000,
11'b10100000110,
11'b10100000111,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b11000000101,
11'b11000000110,
11'b11000000111,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11000100110,
11'b11000100111,
11'b11100000101,
11'b11100000110,
11'b11100000111,
11'b11100010101,
11'b11100010110,
11'b11100010111,
11'b11100100101,
11'b11100100110,
11'b11100100111: edge_mask_reg_512p7[244] <= 1'b1;
 		default: edge_mask_reg_512p7[244] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b10111010,
11'b100111001,
11'b100111010,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100101,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010100,
11'b10010010101,
11'b10010100100,
11'b10010100101,
11'b10101010100,
11'b10101010101,
11'b10101100100,
11'b10101100101,
11'b10101110100,
11'b10101110101,
11'b10110000100,
11'b10110000101,
11'b10110010100,
11'b10110010101,
11'b11001100100,
11'b11001110100,
11'b11010000100,
11'b11010010100: edge_mask_reg_512p7[245] <= 1'b1;
 		default: edge_mask_reg_512p7[245] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1010101,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100101,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110101,
11'b1110110,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110000101,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010000101,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011010,
11'b1010011011,
11'b1100111010,
11'b1100111011,
11'b1101000110,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b10001010101,
11'b10001010110,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101010,
11'b10001101011,
11'b10001110101,
11'b10001110110,
11'b10001110111: edge_mask_reg_512p7[246] <= 1'b1;
 		default: edge_mask_reg_512p7[246] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b10001000101,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10101000100,
11'b10101000101,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11001100101,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101: edge_mask_reg_512p7[247] <= 1'b1;
 		default: edge_mask_reg_512p7[247] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010110,
11'b1110010111,
11'b1110100110,
11'b10001000101,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000100,
11'b10110000101,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11001100101,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11010000101,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101,
11'b11101110100,
11'b11101110101,
11'b11110000100,
11'b11110000101: edge_mask_reg_512p7[248] <= 1'b1;
 		default: edge_mask_reg_512p7[248] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100110,
11'b1110100111,
11'b10001000101,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010011,
11'b10110010100,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11001100101,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101,
11'b11101110100: edge_mask_reg_512p7[249] <= 1'b1;
 		default: edge_mask_reg_512p7[249] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101001001,
11'b1101001010,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10100010111,
11'b10100011000,
11'b10100011001,
11'b10100011010,
11'b10100101000,
11'b10100101001,
11'b10100101010,
11'b11000010111,
11'b11000011000,
11'b11000011001,
11'b11000100111,
11'b11000101000,
11'b11000101001,
11'b11000101010,
11'b11100010111,
11'b11100011000,
11'b11100011001,
11'b11100100111,
11'b11100101000,
11'b11100101001: edge_mask_reg_512p7[250] <= 1'b1;
 		default: edge_mask_reg_512p7[250] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1101110101,
11'b1101110110,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b10010010110,
11'b10010010111,
11'b10010100110,
11'b10010100111,
11'b10010110110,
11'b10010110111,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010111,
11'b10011011000,
11'b10110000110,
11'b10110010110,
11'b10110010111,
11'b10110100110,
11'b10110100111,
11'b10110110110,
11'b10110110111,
11'b10111000110,
11'b10111000111,
11'b10111010110,
11'b10111010111,
11'b11010000110,
11'b11010010110,
11'b11010010111,
11'b11010100110,
11'b11010100111,
11'b11010110110,
11'b11010110111,
11'b11011000110,
11'b11011000111,
11'b11011010110,
11'b11011010111,
11'b11110010110,
11'b11110010111,
11'b11110100110,
11'b11110100111,
11'b11110110110,
11'b11110110111,
11'b11111000110,
11'b11111000111,
11'b11111010111: edge_mask_reg_512p7[251] <= 1'b1;
 		default: edge_mask_reg_512p7[251] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[252] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000101001,
11'b1000101010,
11'b1100011001,
11'b1100011010,
11'b10100000111: edge_mask_reg_512p7[253] <= 1'b1;
 		default: edge_mask_reg_512p7[253] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000010111,
11'b1000100110,
11'b1000100111,
11'b1100010110,
11'b1100010111,
11'b11000000101,
11'b11000000110,
11'b11100000101,
11'b11100000110: edge_mask_reg_512p7[254] <= 1'b1;
 		default: edge_mask_reg_512p7[254] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[255] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[256] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000100111,
11'b10000101000,
11'b10000101001,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001010111,
11'b10001011000,
11'b10100000111,
11'b10100001000,
11'b10100010111,
11'b10100011000,
11'b10100011001,
11'b10100100111,
11'b10100101000,
11'b10100101001,
11'b10100110111,
11'b10100111000,
11'b10101000111,
11'b10101001000,
11'b10101010111,
11'b10101011000,
11'b11000000111,
11'b11000001000,
11'b11000010111,
11'b11000011000,
11'b11000100111,
11'b11000101000,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010111,
11'b11001011000,
11'b11100000111,
11'b11100001000,
11'b11100010111,
11'b11100011000,
11'b11100100111,
11'b11100101000,
11'b11100110111,
11'b11100111000,
11'b11101000111,
11'b11101001000,
11'b11101010111: edge_mask_reg_512p7[257] <= 1'b1;
 		default: edge_mask_reg_512p7[257] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100100,
11'b1100100101,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110111,
11'b1100111000,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10100010100,
11'b10100010101,
11'b10100100100: edge_mask_reg_512p7[258] <= 1'b1;
 		default: edge_mask_reg_512p7[258] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[259] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[260] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[261] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[262] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111100,
11'b110001100,
11'b110011100,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001100,
11'b1010001101,
11'b1010011100,
11'b1010011101,
11'b1010101101,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111000,
11'b1101111001,
11'b1101111100,
11'b1101111101,
11'b1110001100,
11'b1110001101,
11'b1110011101,
11'b1110101101,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10000100111,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10000111010,
11'b10000111101,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001001010,
11'b10001001101,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001011010,
11'b10001011101,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101101,
11'b10001101110,
11'b10100010111,
11'b10100011000,
11'b10100100111,
11'b10100101000,
11'b10100110111,
11'b10100111000,
11'b10101000111,
11'b10101001000,
11'b10101011000: edge_mask_reg_512p7[263] <= 1'b1;
 		default: edge_mask_reg_512p7[263] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[264] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001011,
11'b10011011,
11'b10101011,
11'b10111011,
11'b101111100,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011010,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101001,
11'b1011101010,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10010111100,
11'b10010111101,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011001100,
11'b10011001101,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011100,
11'b10011011101,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101100,
11'b10110110111,
11'b10110111000,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b11011000111,
11'b11011001000,
11'b11011010111,
11'b11011011000: edge_mask_reg_512p7[265] <= 1'b1;
 		default: edge_mask_reg_512p7[265] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011011,
11'b10101011,
11'b10111011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b111001011,
11'b1010011100,
11'b1010011101,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011100,
11'b10011011101,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101100,
11'b10011110111,
11'b10011111000,
11'b10011111001,
11'b10111001000,
11'b10111001001,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b10111111000,
11'b11011000111,
11'b11011001000,
11'b11011010111,
11'b11011011000,
11'b11011100111,
11'b11011101000: edge_mask_reg_512p7[266] <= 1'b1;
 		default: edge_mask_reg_512p7[266] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[267] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111010,
11'b11001001,
11'b11001010,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111001010,
11'b1111010101,
11'b1111010110,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10011100100,
11'b10011100101,
11'b10011110101,
11'b10011110110,
11'b10111100100,
11'b10111100101,
11'b10111110101: edge_mask_reg_512p7[268] <= 1'b1;
 		default: edge_mask_reg_512p7[268] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1101010110,
11'b1101010111,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000111,
11'b1111001000,
11'b10001100100,
11'b10001100101,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10101100100,
11'b10101100101,
11'b10101110100,
11'b10101110101,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110100,
11'b10110110101,
11'b11001100100,
11'b11001100101,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11010110101,
11'b11101100100,
11'b11101110100,
11'b11110000100,
11'b11110010100,
11'b11110100100: edge_mask_reg_512p7[269] <= 1'b1;
 		default: edge_mask_reg_512p7[269] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[270] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[271] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[272] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001010,
11'b111001011,
11'b111011010,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101011,
11'b10011110111,
11'b10011111000,
11'b10011111001,
11'b10011111010,
11'b10111000111,
11'b10111001000,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b10111111001,
11'b11011000111,
11'b11011001000,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100110,
11'b11011100111,
11'b11011101000,
11'b11011110110,
11'b11011110111,
11'b11011111000,
11'b11111010111,
11'b11111100111,
11'b11111110111: edge_mask_reg_512p7[273] <= 1'b1;
 		default: edge_mask_reg_512p7[273] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011011,
11'b101001100,
11'b101011100,
11'b101101100,
11'b101111100,
11'b110001100,
11'b110011100,
11'b110101100,
11'b110111100,
11'b1000111100,
11'b1001001100,
11'b1001001101,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001100,
11'b1010001101,
11'b1010011100,
11'b1010011101,
11'b1010101100,
11'b1010101101,
11'b1010111100,
11'b1010111101,
11'b1011001100,
11'b1100111100,
11'b1100111101,
11'b1101001100,
11'b1101001101,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011100,
11'b1110011101,
11'b1110101100,
11'b1110101101,
11'b1110111100,
11'b1110111101,
11'b1111001101,
11'b10001011010,
11'b10001011011,
11'b10001011100,
11'b10001011101,
11'b10001101010,
11'b10001101011,
11'b10001101100,
11'b10001101101,
11'b10001101110,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10001111101,
11'b10001111110,
11'b10010001011,
11'b10010001100,
11'b10010001101,
11'b10010001110,
11'b10010011011,
11'b10010011100,
11'b10010011101,
11'b10101011010,
11'b10101011011,
11'b10101101001,
11'b10101101010,
11'b10101101011,
11'b10101101100,
11'b10101111001,
11'b10101111010,
11'b10101111011,
11'b10101111100,
11'b10110001010,
11'b10110001011,
11'b10110001100,
11'b10110011011,
11'b10110011100,
11'b11001011010,
11'b11001011011,
11'b11001101001,
11'b11001101010,
11'b11001101011,
11'b11001101100,
11'b11001111001,
11'b11001111010,
11'b11001111011,
11'b11001111100,
11'b11010001001,
11'b11010001010,
11'b11010001011,
11'b11010001100,
11'b11010011011,
11'b11101101001,
11'b11101101010,
11'b11101101011,
11'b11101111001,
11'b11101111010,
11'b11101111011,
11'b11110001001,
11'b11110001010,
11'b11110001011: edge_mask_reg_512p7[274] <= 1'b1;
 		default: edge_mask_reg_512p7[274] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101011,
11'b101001100,
11'b101011100,
11'b101101100,
11'b101111100,
11'b110001100,
11'b110011100,
11'b110101100,
11'b110111100,
11'b1001001100,
11'b1001001101,
11'b1001011100,
11'b1001011101,
11'b1001101100,
11'b1001101101,
11'b1001111100,
11'b1001111101,
11'b1010001100,
11'b1010001101,
11'b1010011100,
11'b1010011101,
11'b1010101100,
11'b1010101101,
11'b1010111100,
11'b1010111101,
11'b1011001100,
11'b1101001100,
11'b1101001101,
11'b1101011100,
11'b1101011101,
11'b1101101100,
11'b1101101101,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001100,
11'b1111001101,
11'b1111011100,
11'b10001101011,
11'b10001101100,
11'b10001101101,
11'b10001101110,
11'b10001111011,
11'b10001111100,
11'b10001111101,
11'b10001111110,
11'b10010001011,
11'b10010001100,
11'b10010001101,
11'b10010001110,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10010011101,
11'b10010011110,
11'b10010101010,
11'b10010101011,
11'b10010101100,
11'b10010101101,
11'b10010111010,
11'b10010111011,
11'b10010111100,
11'b10010111101,
11'b10101101011,
11'b10101101100,
11'b10101111011,
11'b10101111100,
11'b10110001010,
11'b10110001011,
11'b10110001100,
11'b10110011010,
11'b10110011011,
11'b10110011100,
11'b10110101010,
11'b10110101011,
11'b10110101100,
11'b10110111010,
11'b10110111011,
11'b11001101011,
11'b11001101100,
11'b11001111010,
11'b11001111011,
11'b11001111100,
11'b11010001001,
11'b11010001010,
11'b11010001011,
11'b11010001100,
11'b11010011001,
11'b11010011010,
11'b11010011011,
11'b11010011100,
11'b11010101001,
11'b11010101010,
11'b11010101011,
11'b11010111010,
11'b11010111011,
11'b11101101011,
11'b11101111010,
11'b11101111011,
11'b11110001001,
11'b11110001010,
11'b11110001011,
11'b11110011001,
11'b11110011010,
11'b11110011011,
11'b11110101001,
11'b11110101010,
11'b11110101011: edge_mask_reg_512p7[275] <= 1'b1;
 		default: edge_mask_reg_512p7[275] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b1001000110,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110110,
11'b1010110111,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100110,
11'b1110100111,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110101,
11'b10001110110,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010110,
11'b10010010111,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b11001100100,
11'b11001100101,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000100,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010100,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11101100100,
11'b11101100101,
11'b11101110100,
11'b11101110101,
11'b11101110110,
11'b11110000100,
11'b11110000101,
11'b11110000110,
11'b11110000111,
11'b11110010100,
11'b11110010101,
11'b11110010110,
11'b11110010111,
11'b11110100101,
11'b11110100110: edge_mask_reg_512p7[276] <= 1'b1;
 		default: edge_mask_reg_512p7[276] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b1000101010,
11'b1000101011,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b10000011001,
11'b10000011010,
11'b10000011011,
11'b10000101010,
11'b10000101011,
11'b10100001001,
11'b10100011001,
11'b10100011010,
11'b10100101001,
11'b10100101010,
11'b11000001000,
11'b11000001001,
11'b11000001010,
11'b11000011000,
11'b11000011001,
11'b11000011010,
11'b11000101001,
11'b11000101010,
11'b11100001000,
11'b11100001001,
11'b11100001010,
11'b11100011000,
11'b11100011001,
11'b11100011010,
11'b11100101001,
11'b11100101010: edge_mask_reg_512p7[277] <= 1'b1;
 		default: edge_mask_reg_512p7[277] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b100110101,
11'b100110110,
11'b100110111,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110110110,
11'b110110111,
11'b110111000,
11'b1000110101,
11'b1000110110,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b10001000011,
11'b10001010011,
11'b10001010100,
11'b10001100011,
11'b10001100100,
11'b10001110011,
11'b10001110100,
11'b10010000011,
11'b10010000100,
11'b10010010011,
11'b10010100011,
11'b10101010011,
11'b10101100011,
11'b10101110011,
11'b10110000011,
11'b10110010011: edge_mask_reg_512p7[278] <= 1'b1;
 		default: edge_mask_reg_512p7[278] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b100111011,
11'b101001011,
11'b101001100,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b1000101010,
11'b1000101011,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1100011010,
11'b1100011011,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101011,
11'b1101101100,
11'b10000011010,
11'b10000011011,
11'b10000101010,
11'b10000101011,
11'b10000101100,
11'b10000111001,
11'b10000111010,
11'b10000111011,
11'b10000111100,
11'b10000111101,
11'b10001001010,
11'b10001001011,
11'b10100011010,
11'b10100011011,
11'b10100011100,
11'b10100101001,
11'b10100101010,
11'b10100101011,
11'b10100101100,
11'b10100111001,
11'b10100111010,
11'b10100111011,
11'b10101001001,
11'b10101001010,
11'b11000001010,
11'b11000001011,
11'b11000011001,
11'b11000011010,
11'b11000011011,
11'b11000101001,
11'b11000101010,
11'b11000101011,
11'b11000111001,
11'b11000111010,
11'b11000111011,
11'b11001001001,
11'b11001001010,
11'b11100001010,
11'b11100001011,
11'b11100011001,
11'b11100011010,
11'b11100011011,
11'b11100101000,
11'b11100101001,
11'b11100101010,
11'b11100101011,
11'b11100111000,
11'b11100111001,
11'b11100111010,
11'b11101001001,
11'b11101001010: edge_mask_reg_512p7[279] <= 1'b1;
 		default: edge_mask_reg_512p7[279] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010111,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10100010100,
11'b10100010101,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100110011,
11'b10100110100,
11'b10101000011,
11'b10101000100,
11'b11000010100,
11'b11000100100: edge_mask_reg_512p7[280] <= 1'b1;
 		default: edge_mask_reg_512p7[280] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b1000110,
11'b1000111,
11'b1001000,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b101000110,
11'b101000111,
11'b101001000,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1001000110,
11'b1001000111,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110011,
11'b1100110100,
11'b1100110110,
11'b1100110111,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000110011,
11'b10000110100,
11'b10100010100,
11'b10100010101,
11'b10100100011,
11'b10100100100,
11'b10100110011,
11'b11000010100: edge_mask_reg_512p7[281] <= 1'b1;
 		default: edge_mask_reg_512p7[281] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101011000,
11'b1101011001,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10100000110,
11'b10100000111,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10101000111,
11'b10101001000,
11'b11000000101,
11'b11000000110,
11'b11000000111,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11000100110,
11'b11000100111,
11'b11000101000,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000111,
11'b11100000101,
11'b11100000110,
11'b11100000111,
11'b11100010101,
11'b11100010110,
11'b11100010111,
11'b11100100110,
11'b11100100111,
11'b11100110110,
11'b11100110111,
11'b11101000111: edge_mask_reg_512p7[282] <= 1'b1;
 		default: edge_mask_reg_512p7[282] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b100111010,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101001001,
11'b1101001010,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101001,
11'b1110101010,
11'b10001011001,
11'b10001011010,
11'b10001101001,
11'b10001101010,
11'b10001111001,
11'b10001111010,
11'b10010001001,
11'b10010001010,
11'b10101011001,
11'b10101011010,
11'b10101101001,
11'b10101101010,
11'b10101111001,
11'b10101111010,
11'b10110001001,
11'b10110001010,
11'b11001011001,
11'b11001011010,
11'b11001101001,
11'b11001101010,
11'b11001111001,
11'b11001111010,
11'b11010001001,
11'b11010001010,
11'b11010011010,
11'b11101011001,
11'b11101011010,
11'b11101101001,
11'b11101101010,
11'b11101111001,
11'b11101111010,
11'b11110001000,
11'b11110001001,
11'b11110001010: edge_mask_reg_512p7[283] <= 1'b1;
 		default: edge_mask_reg_512p7[283] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011001,
11'b1010011010,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10001001001,
11'b10001001010,
11'b10001001011,
11'b10001011001,
11'b10001011010,
11'b10001011011,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001111001,
11'b10001111010,
11'b10101001001,
11'b10101001010,
11'b10101001011,
11'b10101011001,
11'b10101011010,
11'b10101011011,
11'b10101101001,
11'b10101101010,
11'b10101101011,
11'b10101111001,
11'b10101111010,
11'b11001001001,
11'b11001001010,
11'b11001001011,
11'b11001011001,
11'b11001011010,
11'b11001011011,
11'b11001101001,
11'b11001101010,
11'b11001101011,
11'b11001111001,
11'b11001111010,
11'b11101001010,
11'b11101001011,
11'b11101011001,
11'b11101011010,
11'b11101011011,
11'b11101101001,
11'b11101101010,
11'b11101101011,
11'b11101111001,
11'b11101111010: edge_mask_reg_512p7[284] <= 1'b1;
 		default: edge_mask_reg_512p7[284] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101011,
11'b1111011,
11'b10001011,
11'b10011011,
11'b10101011,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b101111011,
11'b101111100,
11'b110001011,
11'b110001100,
11'b110011100,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b111001011,
11'b1001001100,
11'b1001001101,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001100,
11'b1011011100,
11'b1101001101,
11'b1101011100,
11'b1101011101,
11'b1101101100,
11'b1101101101,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001100,
11'b1111001101,
11'b1111011100,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10010001010,
11'b10010001011,
11'b10010001100,
11'b10010001101,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10010011101,
11'b10010101010,
11'b10010101011,
11'b10010101100,
11'b10010101101,
11'b10010111011,
11'b10010111100,
11'b10010111101,
11'b10011001011,
11'b10011001100,
11'b10011001101,
11'b10101111010,
11'b10101111011,
11'b10110001010,
11'b10110001011,
11'b10110011010,
11'b10110011011,
11'b10110011100,
11'b10110101010,
11'b10110101011,
11'b10110101100,
11'b10110111010,
11'b10110111011,
11'b10110111100,
11'b10111001011,
11'b10111001100,
11'b11001111010,
11'b11001111011,
11'b11010001010,
11'b11010001011,
11'b11010011001,
11'b11010011010,
11'b11010011011,
11'b11010101010,
11'b11010101011,
11'b11010101100,
11'b11010111010,
11'b11010111011,
11'b11010111100,
11'b11011001011,
11'b11011001100,
11'b11110001001,
11'b11110001010,
11'b11110001011,
11'b11110011001,
11'b11110011010,
11'b11110011011,
11'b11110101010,
11'b11110101011,
11'b11110111010,
11'b11110111011,
11'b11111001011: edge_mask_reg_512p7[285] <= 1'b1;
 		default: edge_mask_reg_512p7[285] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[286] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101010,
11'b10101011,
11'b10111010,
11'b10111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b1001001011,
11'b1001001100,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001011,
11'b1011001100,
11'b1101001011,
11'b1101001100,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001100,
11'b10001101010,
11'b10001101011,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010001100,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10101101001,
11'b10101101010,
11'b10101111001,
11'b10101111010,
11'b10101111011,
11'b10110001001,
11'b10110001010,
11'b10110001011,
11'b10110011001,
11'b10110011010,
11'b10110011011,
11'b11001101001,
11'b11001101010,
11'b11001111001,
11'b11001111010,
11'b11010001000,
11'b11010001001,
11'b11010001010,
11'b11010011000,
11'b11010011001,
11'b11010011010,
11'b11101101001,
11'b11101101010,
11'b11101111000,
11'b11101111001,
11'b11101111010,
11'b11110001000,
11'b11110001001,
11'b11110001010,
11'b11110011000,
11'b11110011001,
11'b11110011010: edge_mask_reg_512p7[287] <= 1'b1;
 		default: edge_mask_reg_512p7[287] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[288] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[289] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101010,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101010,
11'b1111101011,
11'b10010011010,
11'b10010101001,
11'b10010101010,
11'b10010101011,
11'b10010111001,
11'b10010111010,
11'b10010111011,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10110011001,
11'b10110011010,
11'b10110101001,
11'b10110101010,
11'b10110111000,
11'b10110111001,
11'b10110111010,
11'b10111001000,
11'b10111001001,
11'b10111001010,
11'b11010011001,
11'b11010011010,
11'b11010101000,
11'b11010101001,
11'b11010101010,
11'b11010111000,
11'b11010111001,
11'b11010111010,
11'b11011001000,
11'b11011001001,
11'b11011001010,
11'b11110011001,
11'b11110101000,
11'b11110101001,
11'b11110101010,
11'b11110111000,
11'b11110111001,
11'b11110111010,
11'b11111001000,
11'b11111001001,
11'b11111001010: edge_mask_reg_512p7[290] <= 1'b1;
 		default: edge_mask_reg_512p7[290] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[291] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100111010,
11'b100111011,
11'b101001011,
11'b101001100,
11'b101011100,
11'b1000011001,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111011,
11'b1000111100,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011100,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111011,
11'b1100111100,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101011100,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10000011011,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000101100,
11'b10100000111,
11'b10100001000,
11'b10100010111,
11'b10100011000,
11'b10100011001,
11'b10100101000,
11'b10100101001,
11'b11000000111,
11'b11000001000,
11'b11000010111,
11'b11000011000,
11'b11000101000,
11'b11100000111,
11'b11100001000,
11'b11100010111,
11'b11100011000: edge_mask_reg_512p7[292] <= 1'b1;
 		default: edge_mask_reg_512p7[292] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000101010,
11'b1000101011,
11'b1000111011,
11'b1000111100,
11'b1100011000,
11'b1100011001,
11'b1100011011,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111011,
11'b1100111100,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10100000111,
11'b10100001000,
11'b10100010111,
11'b10100011000,
11'b10100011001,
11'b11000000111,
11'b11000001000,
11'b11100000111,
11'b11100001000: edge_mask_reg_512p7[293] <= 1'b1;
 		default: edge_mask_reg_512p7[293] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000101010,
11'b1000101011,
11'b1000111011,
11'b1000111100,
11'b1100011000,
11'b1100011001,
11'b1100011011,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111011,
11'b1100111100,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10100000111,
11'b10100001000,
11'b10100011000,
11'b10100011001,
11'b11000000111,
11'b11000001000,
11'b11100000111,
11'b11100001000: edge_mask_reg_512p7[294] <= 1'b1;
 		default: edge_mask_reg_512p7[294] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011101001,
11'b1111101001,
11'b1111101010,
11'b10111110111: edge_mask_reg_512p7[295] <= 1'b1;
 		default: edge_mask_reg_512p7[295] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[296] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b1000110111,
11'b1000111000,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110110,
11'b1110110111,
11'b10001000100,
11'b10001000101,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100100,
11'b10010100101,
11'b10101000100,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b11001010100,
11'b11001100100,
11'b11001100101,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010100100: edge_mask_reg_512p7[297] <= 1'b1;
 		default: edge_mask_reg_512p7[297] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11001000,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1111011000,
11'b1111011001,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011100100: edge_mask_reg_512p7[298] <= 1'b1;
 		default: edge_mask_reg_512p7[298] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101011,
11'b100100110,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101100,
11'b1010101101,
11'b1100100111,
11'b1100101011,
11'b1100101100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b10000111011,
11'b10000111100,
11'b10001001011,
11'b10001001100,
11'b10001010111,
11'b10001011000,
11'b10001011100,
11'b10001100111,
11'b10001101100,
11'b10001111100: edge_mask_reg_512p7[299] <= 1'b1;
 		default: edge_mask_reg_512p7[299] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101010011,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010011,
11'b1110010100,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101001,
11'b1110101010,
11'b10001100011,
11'b10001110011,
11'b10010000011: edge_mask_reg_512p7[300] <= 1'b1;
 		default: edge_mask_reg_512p7[300] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101010011,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101001,
11'b1110101010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010100,
11'b10010010101,
11'b10101110011,
11'b10101110100,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p7[301] <= 1'b1;
 		default: edge_mask_reg_512p7[301] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1101010011,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001001,
11'b1111001010,
11'b10001100011,
11'b10001110011,
11'b10001110100,
11'b10010000011,
11'b10010000100,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110100,
11'b10010110101,
11'b10110000011,
11'b10110000100,
11'b10110010011,
11'b10110010100,
11'b10110100100,
11'b10110110100: edge_mask_reg_512p7[302] <= 1'b1;
 		default: edge_mask_reg_512p7[302] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111000,
11'b10111001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101010011,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100011,
11'b1110101000,
11'b1110101001,
11'b10001100011,
11'b10001110011,
11'b10001110100,
11'b10010000011,
11'b10010000100,
11'b10010010011,
11'b10010010100: edge_mask_reg_512p7[303] <= 1'b1;
 		default: edge_mask_reg_512p7[303] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011001,
11'b1011011010,
11'b1101010011,
11'b1101010100,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111001001,
11'b1111001010,
11'b1111011010,
11'b10001100011,
11'b10001110011,
11'b10010000011,
11'b10010000100,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10011000101,
11'b10110010011,
11'b10110010100,
11'b10110100011,
11'b10110100100,
11'b10110110100: edge_mask_reg_512p7[304] <= 1'b1;
 		default: edge_mask_reg_512p7[304] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001010,
11'b1011001011,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001010,
11'b1111001011,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101010,
11'b10001101011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111010,
11'b10001111011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010001010,
11'b10010001011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011010,
11'b10010011011,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101010,
11'b10101010101,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b10110000111: edge_mask_reg_512p7[305] <= 1'b1;
 		default: edge_mask_reg_512p7[305] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101001,
11'b1011101010,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111010111,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111101001,
11'b1111101010,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011010,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010101010,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10010111010,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10011010110,
11'b10110000101,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10111000101,
11'b10111000110,
11'b11010100101,
11'b11010110101,
11'b11011000101: edge_mask_reg_512p7[306] <= 1'b1;
 		default: edge_mask_reg_512p7[306] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111011,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b101111011,
11'b101111100,
11'b110001100,
11'b1000101010,
11'b1000101011,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001100,
11'b1010001101,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111100,
11'b1101111101,
11'b1110001100,
11'b1110001101,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10000100111,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000101011,
11'b10000101100,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10000111010,
11'b10000111011,
11'b10000111100,
11'b10000111101,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001001010,
11'b10001001011,
11'b10001001100,
11'b10001001101,
11'b10001011000,
11'b10001011001,
11'b10001011010,
11'b10001011011,
11'b10001011100,
11'b10001011101,
11'b10100011000,
11'b10100011001,
11'b10100100111,
11'b10100101000,
11'b10100101001,
11'b10100101010,
11'b10100110111,
11'b10100111000,
11'b10100111001,
11'b10100111010,
11'b10101000111,
11'b10101001000,
11'b10101001001,
11'b10101001010,
11'b10101011000,
11'b10101011001,
11'b10101011010,
11'b11000011000,
11'b11000011001,
11'b11000100111,
11'b11000101000,
11'b11000101001,
11'b11000110111,
11'b11000111000,
11'b11000111001,
11'b11001001000,
11'b11001001001: edge_mask_reg_512p7[307] <= 1'b1;
 		default: edge_mask_reg_512p7[307] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b1000011001,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101011,
11'b1001101100,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000101011,
11'b10000111001,
11'b10000111010,
11'b10000111011,
11'b10001001001,
11'b10001001010,
11'b10100000111,
11'b10100001000,
11'b10100001001,
11'b10100010111,
11'b10100011000,
11'b10100011001,
11'b10100011010,
11'b10100101000,
11'b10100101001,
11'b10100101010,
11'b10100111000,
11'b10100111001,
11'b10100111010,
11'b10101001001,
11'b10101001010,
11'b11000000110,
11'b11000000111,
11'b11000001000,
11'b11000010110,
11'b11000010111,
11'b11000011000,
11'b11000011001,
11'b11000100111,
11'b11000101000,
11'b11000101001,
11'b11000101010,
11'b11000111000,
11'b11000111001,
11'b11000111010,
11'b11001001001,
11'b11001001010,
11'b11100000110,
11'b11100000111,
11'b11100001000,
11'b11100010110,
11'b11100010111,
11'b11100011000,
11'b11100011001,
11'b11100100111,
11'b11100101000,
11'b11100101001,
11'b11100111000,
11'b11100111001,
11'b11100111010,
11'b11101001001: edge_mask_reg_512p7[308] <= 1'b1;
 		default: edge_mask_reg_512p7[308] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011011011,
11'b1011101010,
11'b1111101010,
11'b1111101011,
11'b10111110111,
11'b10111111000: edge_mask_reg_512p7[309] <= 1'b1;
 		default: edge_mask_reg_512p7[309] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101101011,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101010,
11'b1101111010,
11'b1101111011,
11'b1110000110,
11'b1110000111,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b10010000110,
11'b10010000111,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101010,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111010,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110100,
11'b10110110101,
11'b10111000100,
11'b10111000101,
11'b11010010101,
11'b11010100101: edge_mask_reg_512p7[310] <= 1'b1;
 		default: edge_mask_reg_512p7[310] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101010,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010111010,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10110100100,
11'b10110100101,
11'b10110110100,
11'b10110110101,
11'b10111000100,
11'b10111000101: edge_mask_reg_512p7[311] <= 1'b1;
 		default: edge_mask_reg_512p7[311] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111111000,
11'b1111111001,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011010111,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10011110101,
11'b10011110110,
11'b10111000100,
11'b10111000101,
11'b10111000110,
11'b10111010100,
11'b10111010101,
11'b10111010110,
11'b10111100100,
11'b10111100101,
11'b10111100110,
11'b10111110100,
11'b10111110101,
11'b11011000100,
11'b11011000101,
11'b11011010100,
11'b11011010101,
11'b11011100100,
11'b11011100101,
11'b11011110100,
11'b11111010100,
11'b11111100100,
11'b11111110100: edge_mask_reg_512p7[312] <= 1'b1;
 		default: edge_mask_reg_512p7[312] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110001000,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011001000,
11'b10011001001,
11'b10110010111,
11'b10110100111,
11'b10110101000,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b10111001000,
11'b11010010111,
11'b11010100111,
11'b11010101000,
11'b11010110111,
11'b11010111000,
11'b11010111001,
11'b11011000111,
11'b11011001000,
11'b11110100111,
11'b11110101000,
11'b11110110111,
11'b11110111000,
11'b11111000111,
11'b11111001000: edge_mask_reg_512p7[313] <= 1'b1;
 		default: edge_mask_reg_512p7[313] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110001000,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010100111,
11'b10010101000,
11'b10010110111,
11'b10010111000,
11'b10011000111,
11'b10011001000,
11'b10011010111,
11'b10011011000,
11'b10011100111,
11'b10011101000,
11'b10110010111,
11'b10110100111,
11'b10110101000,
11'b10110110111,
11'b10110111000,
11'b10111000111,
11'b10111001000,
11'b10111010111,
11'b10111011000,
11'b10111100111,
11'b10111101000,
11'b11010010111,
11'b11010100111,
11'b11010101000,
11'b11010110111,
11'b11010111000,
11'b11011000111,
11'b11011001000,
11'b11011010111,
11'b11011011000,
11'b11011100111,
11'b11011101000,
11'b11110100111,
11'b11110101000,
11'b11110110111,
11'b11110111000,
11'b11111000111,
11'b11111001000,
11'b11111010111,
11'b11111011000,
11'b11111100111,
11'b11111101000: edge_mask_reg_512p7[314] <= 1'b1;
 		default: edge_mask_reg_512p7[314] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001010,
11'b111001011,
11'b1001011010,
11'b1001011011,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1101011010,
11'b1101011011,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b10001111001,
11'b10001111010,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010101001,
11'b10010101010,
11'b10010101011,
11'b10101111001,
11'b10101111010,
11'b10110001001,
11'b10110001010,
11'b10110001011,
11'b10110011001,
11'b10110011010,
11'b10110011011,
11'b10110101001,
11'b10110101010,
11'b10110101011,
11'b11001111001,
11'b11001111010,
11'b11010001000,
11'b11010001001,
11'b11010001010,
11'b11010011001,
11'b11010011010,
11'b11010011011,
11'b11010101001,
11'b11010101010,
11'b11101111000,
11'b11101111001,
11'b11101111010,
11'b11110001000,
11'b11110001001,
11'b11110001010,
11'b11110011000,
11'b11110011001,
11'b11110011010,
11'b11110101001,
11'b11110101010: edge_mask_reg_512p7[315] <= 1'b1;
 		default: edge_mask_reg_512p7[315] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[316] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011000,
11'b1111011001,
11'b10001111001,
11'b10001111010,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010101000,
11'b10010101001,
11'b10010111000,
11'b10010111001,
11'b10101111001,
11'b10110001000,
11'b10110001001,
11'b10110001010,
11'b10110011000,
11'b10110011001,
11'b10110101000,
11'b10110101001,
11'b10110111000,
11'b10110111001,
11'b11001111001,
11'b11010001000,
11'b11010001001,
11'b11010011000,
11'b11010011001,
11'b11010101000,
11'b11010101001,
11'b11010111000,
11'b11010111001,
11'b11101111001,
11'b11110001000,
11'b11110001001,
11'b11110011000,
11'b11110011001,
11'b11110101000,
11'b11110101001,
11'b11110111000,
11'b11110111001: edge_mask_reg_512p7[317] <= 1'b1;
 		default: edge_mask_reg_512p7[317] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101010,
11'b1101101001,
11'b1101101010,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b11001110101,
11'b11001110110,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110101,
11'b11010110110,
11'b11011000101,
11'b11011000110,
11'b11101110101,
11'b11101110110,
11'b11110000101,
11'b11110000110,
11'b11110010101,
11'b11110010110,
11'b11110100110: edge_mask_reg_512p7[318] <= 1'b1;
 		default: edge_mask_reg_512p7[318] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[319] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1001000111,
11'b1001001000,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010100,
11'b10010010101,
11'b10101010011,
11'b10101010100,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b11001100100,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11010000101,
11'b11101100100,
11'b11101110100: edge_mask_reg_512p7[320] <= 1'b1;
 		default: edge_mask_reg_512p7[320] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1100110111,
11'b1100111000,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110010111,
11'b1110011000,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b11001010100,
11'b11001100100,
11'b11001110100,
11'b11101010100,
11'b11101100100,
11'b11101110100: edge_mask_reg_512p7[321] <= 1'b1;
 		default: edge_mask_reg_512p7[321] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100111001,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10100000110,
11'b10100000111,
11'b10100001000,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b11000000110,
11'b11000000111,
11'b11000001000,
11'b11000010110,
11'b11000010111,
11'b11100000110,
11'b11100000111,
11'b11100010110,
11'b11100010111: edge_mask_reg_512p7[322] <= 1'b1;
 		default: edge_mask_reg_512p7[322] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101001,
11'b101101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101011000,
11'b1101011001,
11'b10000010101,
11'b10000010110,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10100010100,
11'b10100010101,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b11000100100,
11'b11000100101,
11'b11000100110,
11'b11000110100,
11'b11000110101,
11'b11000110110,
11'b11001000101,
11'b11001000110,
11'b11100100100,
11'b11100100101,
11'b11100110100,
11'b11100110101,
11'b11100110110: edge_mask_reg_512p7[323] <= 1'b1;
 		default: edge_mask_reg_512p7[323] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101001,
11'b101101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101011000,
11'b1101011001,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110110,
11'b10000110111,
11'b10001000110,
11'b10001000111,
11'b10100000110,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b11000000101,
11'b11000000110,
11'b11000010101,
11'b11000010110,
11'b11000100101,
11'b11000100110,
11'b11000110101,
11'b11000110110,
11'b11001000101,
11'b11001000110,
11'b11100000101,
11'b11100000110,
11'b11100010101,
11'b11100010110,
11'b11100100101,
11'b11100100110,
11'b11100110101,
11'b11100110110: edge_mask_reg_512p7[324] <= 1'b1;
 		default: edge_mask_reg_512p7[324] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110001010,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1100011000,
11'b1100011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b10000100110,
11'b10000100111,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b11000100101,
11'b11000100110,
11'b11000110101,
11'b11000110110,
11'b11001000101,
11'b11001000110,
11'b11001010101,
11'b11001010110,
11'b11001100110,
11'b11100110101,
11'b11100110110,
11'b11101000101,
11'b11101000110,
11'b11101010101,
11'b11101010110: edge_mask_reg_512p7[325] <= 1'b1;
 		default: edge_mask_reg_512p7[325] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101001,
11'b101101010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101011000,
11'b1101011001,
11'b10000010110,
11'b10000010111,
11'b10000100110,
11'b10000100111,
11'b10000110110,
11'b10000110111,
11'b10001000110,
11'b10001000111,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b11000010101,
11'b11000010110,
11'b11000100101,
11'b11000100110,
11'b11000110101,
11'b11000110110,
11'b11001000101,
11'b11001000110,
11'b11100010101,
11'b11100010110,
11'b11100100101,
11'b11100100110,
11'b11100110101,
11'b11100110110: edge_mask_reg_512p7[326] <= 1'b1;
 		default: edge_mask_reg_512p7[326] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1100011000,
11'b1100011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101111000,
11'b1101111001,
11'b10000100110,
11'b10000100111,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100110,
11'b10001100111,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100110,
11'b10101100111,
11'b11000100101,
11'b11000100110,
11'b11000110101,
11'b11000110110,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100110,
11'b11100110101,
11'b11100110110,
11'b11101000101,
11'b11101000110,
11'b11101010101,
11'b11101010110: edge_mask_reg_512p7[327] <= 1'b1;
 		default: edge_mask_reg_512p7[327] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011011,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1100011000,
11'b1100011001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b10000100110,
11'b10000100111,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110111,
11'b10101111000,
11'b11000100101,
11'b11000100110,
11'b11000110101,
11'b11000110110,
11'b11000110111,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110111,
11'b11001111000,
11'b11100110101,
11'b11100110110,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101010110,
11'b11101010111,
11'b11101011000,
11'b11101100110,
11'b11101100111,
11'b11101101000: edge_mask_reg_512p7[328] <= 1'b1;
 		default: edge_mask_reg_512p7[328] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[329] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[330] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000011000,
11'b1000011001: edge_mask_reg_512p7[331] <= 1'b1;
 		default: edge_mask_reg_512p7[331] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1101111010,
11'b1101111011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b10010001000,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010101011,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10010111011,
11'b10110000111,
11'b10110001000,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b11010000111,
11'b11010010111,
11'b11010011000,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11010110111,
11'b11010111000,
11'b11110010111,
11'b11110011000,
11'b11110100111,
11'b11110101000,
11'b11110110111,
11'b11110111000: edge_mask_reg_512p7[332] <= 1'b1;
 		default: edge_mask_reg_512p7[332] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101101010,
11'b101101011,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101001,
11'b1011101010,
11'b1101111010,
11'b1101111011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10010001000,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10110000111,
11'b10110001000,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b10111001000,
11'b10111001001,
11'b10111011000,
11'b10111011001,
11'b11010000111,
11'b11010010111,
11'b11010011000,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11010110111,
11'b11010111000,
11'b11010111001,
11'b11011001000,
11'b11011001001,
11'b11011011000,
11'b11011011001,
11'b11110010111,
11'b11110011000,
11'b11110100111,
11'b11110101000,
11'b11110110111,
11'b11110111000,
11'b11110111001,
11'b11111000111,
11'b11111001000,
11'b11111001001,
11'b11111011000: edge_mask_reg_512p7[333] <= 1'b1;
 		default: edge_mask_reg_512p7[333] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101101010,
11'b101101011,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101010,
11'b1101111010,
11'b1101111011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101010,
11'b1111101011,
11'b10010001000,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010101011,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10010111011,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10110000111,
11'b10110001000,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110101010,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b10110111010,
11'b10111001000,
11'b10111001001,
11'b10111001010,
11'b10111011001,
11'b10111011010,
11'b11010000111,
11'b11010010111,
11'b11010011000,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11010110111,
11'b11010111000,
11'b11010111001,
11'b11010111010,
11'b11011001000,
11'b11011001001,
11'b11011001010,
11'b11011011000,
11'b11011011001,
11'b11011011010,
11'b11110010111,
11'b11110011000,
11'b11110100111,
11'b11110101000,
11'b11110101001,
11'b11110110111,
11'b11110111000,
11'b11110111001,
11'b11111001000,
11'b11111001001,
11'b11111001010,
11'b11111011000,
11'b11111011001,
11'b11111011010: edge_mask_reg_512p7[334] <= 1'b1;
 		default: edge_mask_reg_512p7[334] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101101010,
11'b101101011,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011010,
11'b1011011011,
11'b1101111010,
11'b1101111011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111011010,
11'b1111011011,
11'b10010001000,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10110000111,
11'b10110001000,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b11010000111,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11110010110,
11'b11110010111,
11'b11110011000,
11'b11110100110,
11'b11110100111,
11'b11110101000: edge_mask_reg_512p7[335] <= 1'b1;
 		default: edge_mask_reg_512p7[335] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[336] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[337] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[338] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[339] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[340] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110100,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000100,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1001110100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000011,
11'b1011000100,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011101000,
11'b1101110011,
11'b1101110100,
11'b1101111000,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000011,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010011,
11'b1111010100,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b10010000011,
11'b10010000100,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100,
11'b10010110011,
11'b10010110100,
11'b10011000011,
11'b10011000100,
11'b10011010011: edge_mask_reg_512p7[341] <= 1'b1;
 		default: edge_mask_reg_512p7[341] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10100110011,
11'b10100110100,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b11001000100,
11'b11001010100,
11'b11001010101: edge_mask_reg_512p7[342] <= 1'b1;
 		default: edge_mask_reg_512p7[342] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[343] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b100101010,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b101111100,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1100011010,
11'b1100011011,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000101011,
11'b10000101100,
11'b10000111000,
11'b10000111001,
11'b10000111010,
11'b10000111011,
11'b10000111100,
11'b10001001000,
11'b10001001001,
11'b10001001010,
11'b10100101000,
11'b10100101001,
11'b10100101010,
11'b10100111000,
11'b10100111001,
11'b10100111010,
11'b10101001000,
11'b10101001001,
11'b11000101000,
11'b11000101001,
11'b11000111000,
11'b11000111001,
11'b11001001000,
11'b11001001001,
11'b11100101000,
11'b11100101001,
11'b11100111000,
11'b11100111001: edge_mask_reg_512p7[344] <= 1'b1;
 		default: edge_mask_reg_512p7[344] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b100101010,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1100011010,
11'b1100011011,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011100,
11'b1110011101,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000101011,
11'b10000111000,
11'b10000111001,
11'b10000111010,
11'b10000111011,
11'b10000111100,
11'b10001001000,
11'b10001001001,
11'b10001001010,
11'b10001001011,
11'b10001001100,
11'b10001011000,
11'b10001011001,
11'b10001011010,
11'b10001011011,
11'b10001011100,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001101100,
11'b10001111001,
11'b10001111010,
11'b10100101000,
11'b10100101001,
11'b10100111000,
11'b10100111001,
11'b10100111010,
11'b10101001000,
11'b10101001001,
11'b10101001010,
11'b10101011000,
11'b10101011001,
11'b10101011010,
11'b10101101000,
11'b10101101001,
11'b10101101010,
11'b10101111001,
11'b11000101000,
11'b11000101001,
11'b11000111000,
11'b11000111001,
11'b11001001000,
11'b11001001001,
11'b11001011000,
11'b11001011001,
11'b11001101000,
11'b11001101001,
11'b11001111001,
11'b11100101000,
11'b11100111000,
11'b11100111001,
11'b11101001000,
11'b11101001001,
11'b11101011000,
11'b11101011001,
11'b11101101000,
11'b11101101001: edge_mask_reg_512p7[345] <= 1'b1;
 		default: edge_mask_reg_512p7[345] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b100101010,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101011,
11'b101101100,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101011,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10000011011,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000101011,
11'b10000111000,
11'b10000111001,
11'b10000111010,
11'b10000111011,
11'b10001001000,
11'b10001001001,
11'b10100001000,
11'b10100001001,
11'b10100010111,
11'b10100011000,
11'b10100011001,
11'b10100100111,
11'b10100101000,
11'b10100101001,
11'b10100111000,
11'b10100111001,
11'b10101001000,
11'b10101001001,
11'b11000001000,
11'b11000010111,
11'b11000011000,
11'b11000011001,
11'b11000100111,
11'b11000101000,
11'b11000101001,
11'b11000111000,
11'b11000111001,
11'b11001001000,
11'b11001001001,
11'b11100010111,
11'b11100011000,
11'b11100100111,
11'b11100101000,
11'b11100111000,
11'b11100111001: edge_mask_reg_512p7[346] <= 1'b1;
 		default: edge_mask_reg_512p7[346] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110001001,
11'b110001010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1100101000,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101111000,
11'b1101111001,
11'b10000110111,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010111,
11'b10001011000,
11'b10001100111,
11'b10001101000,
11'b10100110111,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100111,
11'b10101101000,
11'b11000110111,
11'b11001000110,
11'b11001000111,
11'b11001010110,
11'b11001010111,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11100110111,
11'b11101000110,
11'b11101000111,
11'b11101010110,
11'b11101010111,
11'b11101100110,
11'b11101100111: edge_mask_reg_512p7[347] <= 1'b1;
 		default: edge_mask_reg_512p7[347] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110001001,
11'b110001010,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101111000,
11'b1101111001,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010111,
11'b10001011000,
11'b10001100111,
11'b10001101000,
11'b10100100110,
11'b10100100111,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100111,
11'b10101101000,
11'b11000100110,
11'b11000100111,
11'b11000110110,
11'b11000110111,
11'b11001000110,
11'b11001000111,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11100110101,
11'b11100110110,
11'b11100110111,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101010110,
11'b11101010111,
11'b11101100110,
11'b11101100111: edge_mask_reg_512p7[348] <= 1'b1;
 		default: edge_mask_reg_512p7[348] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1100111000,
11'b1100111001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101001,
11'b1110101010,
11'b10001000111,
11'b10001001000,
11'b10001010111,
11'b10001011000,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10101000111,
11'b10101001000,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100111,
11'b10101101000,
11'b10101110111,
11'b10101111000,
11'b10110000111,
11'b10110001000,
11'b11001000110,
11'b11001000111,
11'b11001010110,
11'b11001010111,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110111,
11'b11001111000,
11'b11010000111,
11'b11010001000,
11'b11010010111,
11'b11101000110,
11'b11101000111,
11'b11101010110,
11'b11101010111,
11'b11101100110,
11'b11101100111,
11'b11101101000,
11'b11101110110,
11'b11101110111,
11'b11101111000,
11'b11110000110,
11'b11110000111,
11'b11110001000: edge_mask_reg_512p7[349] <= 1'b1;
 		default: edge_mask_reg_512p7[349] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1100111000,
11'b1100111001,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b10001000111,
11'b10001001000,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10101000111,
11'b10101001000,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b11001000110,
11'b11001000111,
11'b11001010110,
11'b11001010111,
11'b11001100101,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000101,
11'b11010000110,
11'b11101000110,
11'b11101000111,
11'b11101010110,
11'b11101010111,
11'b11101100101,
11'b11101100110,
11'b11101100111,
11'b11101110100,
11'b11101110101,
11'b11101110110,
11'b11101110111,
11'b11110000101,
11'b11110000110: edge_mask_reg_512p7[350] <= 1'b1;
 		default: edge_mask_reg_512p7[350] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[351] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[352] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10010010110,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11011000101,
11'b11011000110,
11'b11011000111,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100110,
11'b11011100111,
11'b11011101000,
11'b11110100101,
11'b11110110101,
11'b11110110110,
11'b11111000101,
11'b11111000110,
11'b11111000111,
11'b11111010101,
11'b11111010110,
11'b11111010111,
11'b11111011000,
11'b11111100110,
11'b11111100111,
11'b11111101000: edge_mask_reg_512p7[353] <= 1'b1;
 		default: edge_mask_reg_512p7[353] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110001010,
11'b1110001011,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b11010100110,
11'b11010100111,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100111,
11'b11011101000,
11'b11110100110,
11'b11110100111,
11'b11110110110,
11'b11110110111,
11'b11111000110,
11'b11111000111,
11'b11111010110,
11'b11111010111,
11'b11111011000,
11'b11111100110,
11'b11111100111,
11'b11111101000: edge_mask_reg_512p7[354] <= 1'b1;
 		default: edge_mask_reg_512p7[354] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b1111001,
11'b1111010,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10110100110,
11'b10110100111,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100111,
11'b11011101000,
11'b11110100101,
11'b11110100110,
11'b11110110101,
11'b11110110110,
11'b11111000101,
11'b11111000110,
11'b11111000111,
11'b11111010110,
11'b11111010111,
11'b11111011000,
11'b11111100110,
11'b11111100111,
11'b11111101000: edge_mask_reg_512p7[355] <= 1'b1;
 		default: edge_mask_reg_512p7[355] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001111011,
11'b1001111100,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101001,
11'b1011101010,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10010011000,
11'b10010011001,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010101011,
11'b10010101100,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10010111011,
11'b10010111100,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011100111,
11'b10011101000,
11'b10110011000,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100111,
11'b10111101000,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11010110111,
11'b11010111000,
11'b11010111001,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011001001,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100111,
11'b11011101000,
11'b11110100111,
11'b11110101000,
11'b11110110111,
11'b11110111000,
11'b11111000110,
11'b11111000111,
11'b11111001000,
11'b11111010110,
11'b11111010111: edge_mask_reg_512p7[356] <= 1'b1;
 		default: edge_mask_reg_512p7[356] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110101011,
11'b1110101100,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011011100,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10011101100,
11'b10111000111,
11'b10111001000,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b11011000110,
11'b11011000111,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100110,
11'b11011100111,
11'b11011101000,
11'b11111000110,
11'b11111000111,
11'b11111010110,
11'b11111010111: edge_mask_reg_512p7[357] <= 1'b1;
 		default: edge_mask_reg_512p7[357] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101010,
11'b10101011,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1100111010,
11'b1100111011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110000111,
11'b1110001000,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011010,
11'b10001011011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101010,
11'b10001101011,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111010,
11'b10001111011,
11'b10010000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110101,
11'b10101110110,
11'b10101110111: edge_mask_reg_512p7[358] <= 1'b1;
 		default: edge_mask_reg_512p7[358] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1100011010,
11'b1100011011,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001010,
11'b1110001011,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10000111011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001001011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011010,
11'b10001011011,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101011,
11'b10100100101,
11'b10100110101,
11'b10101000101: edge_mask_reg_512p7[359] <= 1'b1;
 		default: edge_mask_reg_512p7[359] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b1000101011,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1100110100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011010,
11'b10001011011,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101011: edge_mask_reg_512p7[360] <= 1'b1;
 		default: edge_mask_reg_512p7[360] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[361] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110101,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100110,
11'b101100111,
11'b101101000,
11'b1000010111,
11'b1000011000,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101010100,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b10000010100,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001010011,
11'b10001010100,
11'b10100010100,
11'b10100100011,
11'b10100100100,
11'b10100110011,
11'b10100110100,
11'b10101000011,
11'b10101000100,
11'b10101010011,
11'b10101010100: edge_mask_reg_512p7[362] <= 1'b1;
 		default: edge_mask_reg_512p7[362] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011010,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111101001,
11'b10010001001,
11'b10010001010,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10010111000,
11'b10010111001,
11'b10010111010,
11'b10011001000,
11'b10011001001,
11'b10110001001,
11'b10110001010,
11'b10110011000,
11'b10110011001,
11'b10110011010,
11'b10110101000,
11'b10110101001,
11'b10110101010,
11'b10110111000,
11'b10110111001,
11'b10111001000,
11'b10111001001,
11'b11010001001,
11'b11010011000,
11'b11010011001,
11'b11010011010,
11'b11010101000,
11'b11010101001,
11'b11010101010,
11'b11010111000,
11'b11010111001,
11'b11011001000,
11'b11011001001,
11'b11110001001,
11'b11110011000,
11'b11110011001,
11'b11110101000,
11'b11110101001,
11'b11110111000,
11'b11110111001,
11'b11111001000,
11'b11111001001: edge_mask_reg_512p7[363] <= 1'b1;
 		default: edge_mask_reg_512p7[363] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10110100111,
11'b10110101000,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b11010100111,
11'b11010101000,
11'b11010110111,
11'b11010111000,
11'b11010111001,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100110,
11'b11011100111,
11'b11110100111,
11'b11110101000,
11'b11110110111,
11'b11110111000,
11'b11111000110,
11'b11111000111,
11'b11111001000,
11'b11111010110,
11'b11111010111,
11'b11111011000,
11'b11111100101,
11'b11111100110,
11'b11111100111: edge_mask_reg_512p7[364] <= 1'b1;
 		default: edge_mask_reg_512p7[364] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110101000,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10110110110,
11'b10111000110,
11'b10111000111,
11'b10111010110,
11'b10111010111,
11'b10111100110,
11'b10111100111,
11'b11011000110,
11'b11011000111,
11'b11011010110,
11'b11011010111,
11'b11011100110,
11'b11011100111,
11'b11111000110,
11'b11111000111,
11'b11111010101,
11'b11111010110,
11'b11111010111,
11'b11111100101,
11'b11111100110,
11'b11111100111: edge_mask_reg_512p7[365] <= 1'b1;
 		default: edge_mask_reg_512p7[365] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10101001,
11'b10101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000110,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000101,
11'b10010000110,
11'b10101000110,
11'b10101000111,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000101,
11'b10110000110,
11'b11001000110,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11001110110: edge_mask_reg_512p7[366] <= 1'b1;
 		default: edge_mask_reg_512p7[366] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10001010101,
11'b10001010110,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110100,
11'b10010110101,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110110100,
11'b11001100100,
11'b11001100101,
11'b11001110100,
11'b11001110101,
11'b11010000100: edge_mask_reg_512p7[367] <= 1'b1;
 		default: edge_mask_reg_512p7[367] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101011,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011100,
11'b101101100,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011100,
11'b1001011101,
11'b1001101100,
11'b1001101101,
11'b1001111100,
11'b1001111101,
11'b1010001101,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101011100,
11'b1101011101,
11'b1101101100,
11'b1101101101,
11'b1101111101,
11'b1110001101,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000100111,
11'b10000101000,
11'b10000101001,
11'b10000101100,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10000111100,
11'b10000111101,
11'b10001001000,
11'b10001001001,
11'b10001001101,
11'b10100100111,
11'b10100101000,
11'b10100110111,
11'b10100111000: edge_mask_reg_512p7[368] <= 1'b1;
 		default: edge_mask_reg_512p7[368] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1100110100,
11'b1100110101,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011010,
11'b10000110100,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11001110110: edge_mask_reg_512p7[369] <= 1'b1;
 		default: edge_mask_reg_512p7[369] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b100111010,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111010,
11'b1010111011,
11'b1101001001,
11'b1101001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010001010,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b11001100101,
11'b11001100110,
11'b11001110101,
11'b11001110110,
11'b11010000101,
11'b11010000110: edge_mask_reg_512p7[370] <= 1'b1;
 		default: edge_mask_reg_512p7[370] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b100111010,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100110,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010111001,
11'b1010111010,
11'b1101001001,
11'b1101001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100101,
11'b1110100110,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111001,
11'b1110111010,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10101010110,
11'b10101010111,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000100,
11'b11010000101: edge_mask_reg_512p7[371] <= 1'b1;
 		default: edge_mask_reg_512p7[371] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1100111001,
11'b1100111010,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001001,
11'b1110001010,
11'b1110011010,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110101,
11'b11001110110: edge_mask_reg_512p7[372] <= 1'b1;
 		default: edge_mask_reg_512p7[372] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b100111010,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001001,
11'b111001010,
11'b111001011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1101001001,
11'b1101001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110110110,
11'b1110110111,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110110,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100101,
11'b10110100110,
11'b11001100101,
11'b11001100110,
11'b11001110101,
11'b11001110110,
11'b11010000101,
11'b11010000110,
11'b11010010101,
11'b11010100101: edge_mask_reg_512p7[373] <= 1'b1;
 		default: edge_mask_reg_512p7[373] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001010,
11'b100111010,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101001001,
11'b1101001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10101010110,
11'b10101010111,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100101,
11'b10110100110,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101: edge_mask_reg_512p7[374] <= 1'b1;
 		default: edge_mask_reg_512p7[374] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11001000,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1111011000,
11'b1111011001,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011100100: edge_mask_reg_512p7[375] <= 1'b1;
 		default: edge_mask_reg_512p7[375] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[376] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101101010,
11'b101101011,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011010,
11'b1111011011,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101010,
11'b10010101011,
11'b10010110011,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111011,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110101: edge_mask_reg_512p7[377] <= 1'b1;
 		default: edge_mask_reg_512p7[377] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001001,
11'b111001010,
11'b111001011,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001010,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010011010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110011,
11'b10010110100,
11'b10110000100,
11'b10110010100: edge_mask_reg_512p7[378] <= 1'b1;
 		default: edge_mask_reg_512p7[378] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001001,
11'b111001010,
11'b111001011,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1101010101,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001010,
11'b10001010101,
11'b10001100100,
11'b10001100101,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010011010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110011,
11'b10010110100,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010100: edge_mask_reg_512p7[379] <= 1'b1;
 		default: edge_mask_reg_512p7[379] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001001,
11'b111001010,
11'b111001011,
11'b1001011011,
11'b1001100100,
11'b1001100101,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001010,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010011010,
11'b10010100011,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110011,
11'b10010110100: edge_mask_reg_512p7[380] <= 1'b1;
 		default: edge_mask_reg_512p7[380] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000011000,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010110,
11'b10001010111,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b11000110110,
11'b11000110111,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11100110110,
11'b11100110111,
11'b11100111000,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101001000,
11'b11101010101,
11'b11101010110,
11'b11101010111: edge_mask_reg_512p7[381] <= 1'b1;
 		default: edge_mask_reg_512p7[381] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b1000010111,
11'b1000011000,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010110,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010110,
11'b11000110101,
11'b11000110110,
11'b11000110111,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010110,
11'b11100110101,
11'b11100110110,
11'b11100110111,
11'b11100111000,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101001000,
11'b11101010110: edge_mask_reg_512p7[382] <= 1'b1;
 		default: edge_mask_reg_512p7[382] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011001000,
11'b1011001001,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10001100110,
11'b10001100111,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10101100110,
11'b10101100111,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b11001100110,
11'b11001100111,
11'b11001110110,
11'b11001110111,
11'b11010000110,
11'b11010000111,
11'b11010001000,
11'b11010010111,
11'b11010011000,
11'b11010100111,
11'b11010101000,
11'b11101100101,
11'b11101100110,
11'b11101100111,
11'b11101110101,
11'b11101110110,
11'b11101110111,
11'b11110000101,
11'b11110000110,
11'b11110000111,
11'b11110001000,
11'b11110010110,
11'b11110010111,
11'b11110011000,
11'b11110100110,
11'b11110100111,
11'b11110101000: edge_mask_reg_512p7[383] <= 1'b1;
 		default: edge_mask_reg_512p7[383] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10001101000,
11'b10001101001,
11'b10001111000,
11'b10001111001,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010101000,
11'b10010101001,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110101000,
11'b10110101001,
11'b11001101000,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11010000111,
11'b11010001000,
11'b11010001001,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010100111,
11'b11010101000,
11'b11010101001,
11'b11101101000,
11'b11101110111,
11'b11101111000,
11'b11101111001,
11'b11110000111,
11'b11110001000,
11'b11110001001,
11'b11110010111,
11'b11110011000,
11'b11110100111,
11'b11110101000: edge_mask_reg_512p7[384] <= 1'b1;
 		default: edge_mask_reg_512p7[384] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[385] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[386] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[387] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10110010100,
11'b10110010101,
11'b10110100100,
11'b10110100101,
11'b10110110100,
11'b10110110101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11010110101,
11'b11110010100,
11'b11110100100: edge_mask_reg_512p7[388] <= 1'b1;
 		default: edge_mask_reg_512p7[388] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101010101,
11'b101010110,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000110,
11'b1111000111,
11'b10001110100,
11'b10001110101,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110100,
11'b10010110101,
11'b10101110100,
11'b10101110101,
11'b10110000100,
11'b10110000101,
11'b10110010100,
11'b10110010101,
11'b10110100100,
11'b10110100101,
11'b10110110100,
11'b10110110101,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11101110100,
11'b11110000100,
11'b11110010100,
11'b11110100100: edge_mask_reg_512p7[389] <= 1'b1;
 		default: edge_mask_reg_512p7[389] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10110010100,
11'b10110010101,
11'b10110100100,
11'b10110100101,
11'b10110110100,
11'b10110110101,
11'b10111000100,
11'b10111000101,
11'b10111010100,
11'b10111010101,
11'b10111100100,
11'b10111100101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11010110101,
11'b11011000100,
11'b11011000101,
11'b11011010100,
11'b11011010101,
11'b11011100100,
11'b11011100101,
11'b11110010100,
11'b11110100100,
11'b11110110100,
11'b11111000100,
11'b11111010100: edge_mask_reg_512p7[390] <= 1'b1;
 		default: edge_mask_reg_512p7[390] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000101,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1010101,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1110101,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1101010110,
11'b1101010111,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000110,
11'b1111000111,
11'b10001100100,
11'b10001100101,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110100,
11'b10010110101,
11'b10101100100,
11'b10101100101,
11'b10101110100,
11'b10101110101,
11'b10110000100,
11'b10110000101,
11'b10110010100,
11'b10110010101,
11'b10110100100,
11'b10110100101,
11'b10110110100,
11'b10110110101,
11'b11001100100,
11'b11001100101,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11101100100,
11'b11101110100,
11'b11110000100,
11'b11110010100,
11'b11110100100: edge_mask_reg_512p7[391] <= 1'b1;
 		default: edge_mask_reg_512p7[391] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010010110,
11'b1010010111,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b10010110101,
11'b10010110110,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10011010101,
11'b10011010110,
11'b10011010111,
11'b10110110101,
11'b10110110110,
11'b10111000101,
11'b10111000110,
11'b10111010101,
11'b10111010110,
11'b11010110101,
11'b11010110110,
11'b11011000101,
11'b11011000110,
11'b11011010101,
11'b11011010110,
11'b11110110101,
11'b11110110110,
11'b11111000101,
11'b11111000110,
11'b11111010101,
11'b11111010110: edge_mask_reg_512p7[392] <= 1'b1;
 		default: edge_mask_reg_512p7[392] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b10000101,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b101110110,
11'b101110111,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100111,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110101,
11'b10010110110,
11'b10011000101,
11'b10011000110,
11'b10011010101,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10111000101,
11'b10111000110,
11'b10111010101,
11'b11010010100,
11'b11010010101,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11011000101,
11'b11011000110,
11'b11110010101,
11'b11110100100,
11'b11110100101,
11'b11110110100,
11'b11110110101,
11'b11110110110,
11'b11111000100,
11'b11111000101,
11'b11111000110: edge_mask_reg_512p7[393] <= 1'b1;
 		default: edge_mask_reg_512p7[393] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1110000111,
11'b1110001000,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111100111,
11'b10010010101,
11'b10010010110,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10011000101,
11'b10011000110,
11'b10011010101,
11'b10110010101,
11'b10110010110,
11'b10110100101,
11'b10110100110,
11'b10110110101,
11'b10110110110,
11'b10111000101,
11'b10111000110,
11'b10111010101,
11'b11010010101,
11'b11010010110,
11'b11010100101,
11'b11010100110,
11'b11010110101,
11'b11010110110,
11'b11011000101,
11'b11011000110,
11'b11110010101,
11'b11110100100,
11'b11110100101,
11'b11110100110,
11'b11110110101,
11'b11110110110,
11'b11111000101,
11'b11111000110: edge_mask_reg_512p7[394] <= 1'b1;
 		default: edge_mask_reg_512p7[394] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[395] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111001,
11'b10111010,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111010,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111001001,
11'b1111001010,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111001,
11'b10011010101,
11'b10011010110,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10011110101,
11'b10011110110,
11'b10011110111,
11'b10111100100,
11'b10111100101,
11'b10111100110,
11'b10111110100,
11'b10111110101,
11'b10111110110,
11'b11011100100,
11'b11011100101,
11'b11011110100,
11'b11011110101: edge_mask_reg_512p7[396] <= 1'b1;
 		default: edge_mask_reg_512p7[396] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111001,
11'b10111010,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111010,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111001001,
11'b1111001010,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011110101,
11'b10011110110,
11'b10111100011,
11'b10111100100,
11'b10111100101,
11'b10111110100,
11'b10111110101,
11'b11011100100,
11'b11011110100: edge_mask_reg_512p7[397] <= 1'b1;
 		default: edge_mask_reg_512p7[397] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[398] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101101001,
11'b1101101010,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b10101010110,
11'b11000100100,
11'b11000100101,
11'b11000100110,
11'b11000110100,
11'b11000110101,
11'b11000110110,
11'b11001000101,
11'b11001000110,
11'b11100100100,
11'b11100100101,
11'b11100110100,
11'b11100110101,
11'b11101000101: edge_mask_reg_512p7[399] <= 1'b1;
 		default: edge_mask_reg_512p7[399] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1100011001,
11'b1100011010,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b10000100111,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110101,
11'b10101110110,
11'b11000110101,
11'b11000110110,
11'b11001000101,
11'b11001000110,
11'b11001010101,
11'b11001010110,
11'b11001100101,
11'b11001100110,
11'b11001110101,
11'b11001110110,
11'b11100110101,
11'b11101000101,
11'b11101010101,
11'b11101010110,
11'b11101100101,
11'b11101100110,
11'b11101110101,
11'b11101110110: edge_mask_reg_512p7[400] <= 1'b1;
 		default: edge_mask_reg_512p7[400] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101011010,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10100000110,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100110110,
11'b10100110111,
11'b11000000101,
11'b11000010100,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11000100101,
11'b11000100110,
11'b11000100111,
11'b11000110110,
11'b11000110111,
11'b11100010101,
11'b11100010110,
11'b11100100101,
11'b11100100110,
11'b11100110110: edge_mask_reg_512p7[401] <= 1'b1;
 		default: edge_mask_reg_512p7[401] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101011000,
11'b1101011001,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100110101,
11'b10100110110,
11'b10101000101,
11'b10101000110,
11'b11000000101,
11'b11000010100,
11'b11000010101,
11'b11000010110,
11'b11000100100,
11'b11000100101,
11'b11000100110,
11'b11000110100,
11'b11000110101,
11'b11000110110,
11'b11100010100,
11'b11100010101,
11'b11100100100,
11'b11100100101,
11'b11100110100,
11'b11100110101: edge_mask_reg_512p7[402] <= 1'b1;
 		default: edge_mask_reg_512p7[402] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011010,
11'b1011011,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011010,
11'b10011011,
11'b10101010,
11'b10101011,
11'b10111010,
11'b10111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001011,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001011,
11'b1011001100,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001011,
11'b1111001100,
11'b1111001101,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010001100,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10010101000,
11'b10010101001,
11'b10010101010,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110001010,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110011010,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110101010,
11'b11001100111,
11'b11001101000,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11010000111,
11'b11010001000,
11'b11010001001,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010100111,
11'b11010101000,
11'b11010101001: edge_mask_reg_512p7[403] <= 1'b1;
 		default: edge_mask_reg_512p7[403] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111010,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100101,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b11001100111,
11'b11001101000,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11010000111,
11'b11010001000: edge_mask_reg_512p7[404] <= 1'b1;
 		default: edge_mask_reg_512p7[404] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011011,
11'b1101011,
11'b1111011,
11'b10001011,
11'b10011011,
11'b10101011,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b1000101000,
11'b1000101011,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1100101011,
11'b1100101100,
11'b1100110111,
11'b1100111000,
11'b1100111011,
11'b1100111100,
11'b1100111101,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001011,
11'b1101001100,
11'b1101001101,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011011,
11'b1101011100,
11'b1101011101,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101110111,
11'b1101111000,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110000111,
11'b1110001000,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101100,
11'b1110101101,
11'b10001001100,
11'b10001001101,
11'b10001011100,
11'b10001011101,
11'b10001101100,
11'b10001101101,
11'b10001111100,
11'b10001111101: edge_mask_reg_512p7[405] <= 1'b1;
 		default: edge_mask_reg_512p7[405] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111011000,
11'b1111011001,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10011000101,
11'b10011000110,
11'b10110010101,
11'b10110010110,
11'b10110100101,
11'b10110100110,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10111000101,
11'b11010010101,
11'b11010010110,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010110100,
11'b11010110101,
11'b11110100101,
11'b11110110101: edge_mask_reg_512p7[406] <= 1'b1;
 		default: edge_mask_reg_512p7[406] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111000,
11'b1111001,
11'b1111010,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101001,
11'b1011101010,
11'b1110010101,
11'b1110010110,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b10010010101,
11'b10010010110,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000101,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10110010101,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b11010100100,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110100,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11110100101,
11'b11110100110,
11'b11110110101,
11'b11110110110,
11'b11110110111: edge_mask_reg_512p7[407] <= 1'b1;
 		default: edge_mask_reg_512p7[407] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001101,
11'b1001011101,
11'b1001101101,
11'b1001111101,
11'b1010001101,
11'b1010011101,
11'b1010101101,
11'b1010111101,
11'b1101001101,
11'b1101011101,
11'b1101101101,
11'b1101111100,
11'b1101111101,
11'b1110001100,
11'b1110001101,
11'b1110011100,
11'b1110011101,
11'b1110101100,
11'b1110101101,
11'b1110111100,
11'b1110111101,
11'b1111001101,
11'b10001111011,
11'b10001111100,
11'b10001111101,
11'b10001111110,
11'b10010001011,
11'b10010001100,
11'b10010001101,
11'b10010001110,
11'b10010011011,
11'b10010011100,
11'b10010011101,
11'b10010011110,
11'b10010101011,
11'b10010101100,
11'b10010101101,
11'b10010101110,
11'b10010111100,
11'b10010111101,
11'b10011001101,
11'b10101111011,
11'b10101111100,
11'b10101111101,
11'b10110001011,
11'b10110001100,
11'b10110001101,
11'b10110011011,
11'b10110011100,
11'b10110011101,
11'b10110101011,
11'b10110101100,
11'b10110101101,
11'b10110111100,
11'b10110111101,
11'b10111001101,
11'b11001111011,
11'b11001111100,
11'b11010001010,
11'b11010001011,
11'b11010001100,
11'b11010001101,
11'b11010011011,
11'b11010011100,
11'b11010011101,
11'b11010101011,
11'b11010101100,
11'b11010101101,
11'b11010111100,
11'b11010111101,
11'b11101111011,
11'b11110001010,
11'b11110001011,
11'b11110001100,
11'b11110011010,
11'b11110011011,
11'b11110011100,
11'b11110101011,
11'b11110101100,
11'b11110111100: edge_mask_reg_512p7[408] <= 1'b1;
 		default: edge_mask_reg_512p7[408] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100101000,
11'b100101001,
11'b100101010,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b10000011000,
11'b10000011001,
11'b10100001000,
11'b10100001001,
11'b10100011000,
11'b10100011001,
11'b11000000111,
11'b11000001000,
11'b11000001001,
11'b11000011000,
11'b11000011001,
11'b11100000111,
11'b11100001000,
11'b11100001001,
11'b11100011000: edge_mask_reg_512p7[409] <= 1'b1;
 		default: edge_mask_reg_512p7[409] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[410] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000111,
11'b1010001000,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b10000100111,
11'b10000101000,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10100100111,
11'b10100101000,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b11000100111,
11'b11000101000,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11001100101,
11'b11001100110,
11'b11100100111,
11'b11100110110,
11'b11100110111,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101010101,
11'b11101010110,
11'b11101010111,
11'b11101100101,
11'b11101100110: edge_mask_reg_512p7[411] <= 1'b1;
 		default: edge_mask_reg_512p7[411] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100101010,
11'b1000011001,
11'b1000101001,
11'b1000101010,
11'b1100011001,
11'b1100011010,
11'b1100101001,
11'b1100101010,
11'b10100001000,
11'b10100001001,
11'b10100011001,
11'b11000001000,
11'b11000001001,
11'b11000011001,
11'b11100001000,
11'b11100001001,
11'b11100011001: edge_mask_reg_512p7[412] <= 1'b1;
 		default: edge_mask_reg_512p7[412] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100101010,
11'b1000011001,
11'b1000101001,
11'b1000101010,
11'b1100011001,
11'b1100011010,
11'b1100101001,
11'b1100101010,
11'b10100001000,
11'b10100001001,
11'b10100011001,
11'b11000001000,
11'b11000001001,
11'b11000011001,
11'b11100001000,
11'b11100001001,
11'b11100011001: edge_mask_reg_512p7[413] <= 1'b1;
 		default: edge_mask_reg_512p7[413] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[414] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[415] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011001,
11'b1110011010,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10100110110,
11'b10100110111,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101011001,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b11000110111,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010110,
11'b11001010111,
11'b11001011000,
11'b11001100111,
11'b11001101000,
11'b11001110111,
11'b11001111000,
11'b11101000110,
11'b11101000111,
11'b11101001000,
11'b11101010110,
11'b11101010111,
11'b11101011000,
11'b11101100110,
11'b11101100111,
11'b11101101000,
11'b11101110110,
11'b11101110111,
11'b11101111000: edge_mask_reg_512p7[416] <= 1'b1;
 		default: edge_mask_reg_512p7[416] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110010110,
11'b110010111,
11'b110011000,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010110,
11'b1010010111,
11'b1100010111,
11'b1100011000,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b10000100101,
11'b10000100110,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10100100100,
11'b10100100101,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101110011,
11'b10101110100,
11'b11000110100,
11'b11000110101,
11'b11000110110,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010100,
11'b11001010101,
11'b11001100100,
11'b11100110100,
11'b11100110101,
11'b11101000100,
11'b11101000101,
11'b11101010100: edge_mask_reg_512p7[417] <= 1'b1;
 		default: edge_mask_reg_512p7[417] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[418] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b10011100110,
11'b10011100111,
11'b10011110101,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111110110,
11'b10111110111: edge_mask_reg_512p7[419] <= 1'b1;
 		default: edge_mask_reg_512p7[419] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[420] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011001,
11'b1001011010,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011010,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000110111,
11'b10000111000,
11'b10100000110,
11'b10100000111,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100110110,
11'b10100110111,
11'b11000000101,
11'b11000000110,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11000100101,
11'b11000100110,
11'b11000100111,
11'b11000110110,
11'b11000110111,
11'b11100000110,
11'b11100010101,
11'b11100010110,
11'b11100100101,
11'b11100100110,
11'b11100110110: edge_mask_reg_512p7[421] <= 1'b1;
 		default: edge_mask_reg_512p7[421] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110111,
11'b101111000,
11'b101111001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110111,
11'b1001111000,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10100110101,
11'b10100110110,
11'b10101000101,
11'b10101000110,
11'b10101010101,
11'b10101010110,
11'b11000110101,
11'b11000110110,
11'b11001000101,
11'b11001000110,
11'b11001010101,
11'b11001010110,
11'b11100110101,
11'b11101000100,
11'b11101000101,
11'b11101000110,
11'b11101010101,
11'b11101010110: edge_mask_reg_512p7[422] <= 1'b1;
 		default: edge_mask_reg_512p7[422] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010010110,
11'b1010010111,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001110101,
11'b10001110110,
11'b10100110101,
11'b10100110110,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b11000110101,
11'b11000110110,
11'b11001000100,
11'b11001000101,
11'b11001000110,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11100110101,
11'b11101000100,
11'b11101000101,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101,
11'b11101110100,
11'b11101110101: edge_mask_reg_512p7[423] <= 1'b1;
 		default: edge_mask_reg_512p7[423] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101111001,
11'b101111010,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001001000,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b11000110101,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000101,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010101,
11'b11001010110,
11'b11001010111,
11'b11100110101,
11'b11100110110,
11'b11100110111,
11'b11101000100,
11'b11101000101,
11'b11101000110,
11'b11101000111,
11'b11101001000,
11'b11101010110,
11'b11101010111: edge_mask_reg_512p7[424] <= 1'b1;
 		default: edge_mask_reg_512p7[424] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[425] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b11000000101,
11'b11000000110,
11'b11000010100,
11'b11000010101,
11'b11100000101,
11'b11100010101: edge_mask_reg_512p7[426] <= 1'b1;
 		default: edge_mask_reg_512p7[426] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011010,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111000110,
11'b10111000111,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b11011000110,
11'b11011000111,
11'b11011010110,
11'b11011010111,
11'b11011100110,
11'b11011100111,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111010110,
11'b11111010111,
11'b11111100110,
11'b11111100111,
11'b11111110101,
11'b11111110110,
11'b11111110111: edge_mask_reg_512p7[427] <= 1'b1;
 		default: edge_mask_reg_512p7[427] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10111000,
11'b10111001,
11'b10111010,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110111001,
11'b110111010,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111010110,
11'b10111010111,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b11011010110,
11'b11011100110,
11'b11011100111,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111100110,
11'b11111100111,
11'b11111110101,
11'b11111110110: edge_mask_reg_512p7[428] <= 1'b1;
 		default: edge_mask_reg_512p7[428] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011010110,
11'b10011010111,
11'b10011100110,
11'b10011100111,
11'b10011110110,
11'b10011110111,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b11011010101,
11'b11011010110,
11'b11011100101,
11'b11011100110,
11'b11011110101,
11'b11011110110,
11'b11111010101,
11'b11111010110,
11'b11111100101,
11'b11111100110,
11'b11111110101,
11'b11111110110: edge_mask_reg_512p7[429] <= 1'b1;
 		default: edge_mask_reg_512p7[429] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111010,
11'b10111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b1001001011,
11'b1001001100,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111011,
11'b1010111100,
11'b1010111101,
11'b1011001011,
11'b1011001100,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110101101,
11'b1110111011,
11'b1110111100,
11'b1110111101,
11'b1111001100,
11'b10001101001,
11'b10001101010,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10001111100,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010001100,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10101101001,
11'b10101111000,
11'b10101111001,
11'b10101111010,
11'b10110001000,
11'b10110001001,
11'b10110001010,
11'b10110011001,
11'b10110011010,
11'b11001101000,
11'b11001101001,
11'b11001111000,
11'b11001111001,
11'b11001111010,
11'b11010001000,
11'b11010001001,
11'b11010001010,
11'b11010011000,
11'b11010011001,
11'b11010011010,
11'b11101111000,
11'b11101111001,
11'b11110001000,
11'b11110001001,
11'b11110011000,
11'b11110011001: edge_mask_reg_512p7[430] <= 1'b1;
 		default: edge_mask_reg_512p7[430] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111010,
11'b1111011,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111011,
11'b110111100,
11'b1001001011,
11'b1001001100,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1001111101,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1101001011,
11'b1101001100,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101101101,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10101101001,
11'b10101101010,
11'b10101111000,
11'b10101111001,
11'b10101111010,
11'b10101111011,
11'b10110001000,
11'b10110001001,
11'b10110001010,
11'b10110001011,
11'b11001101000,
11'b11001101001,
11'b11001101010,
11'b11001111000,
11'b11001111001,
11'b11001111010,
11'b11010001000,
11'b11010001001,
11'b11010001010,
11'b11101101001,
11'b11101101010,
11'b11101111000,
11'b11101111001,
11'b11101111010,
11'b11110001000,
11'b11110001001,
11'b11110001010: edge_mask_reg_512p7[431] <= 1'b1;
 		default: edge_mask_reg_512p7[431] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110101000,
11'b1110101001,
11'b10001000101,
11'b10001000110,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010110,
11'b10010010111,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101100111,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110010110,
11'b10110010111,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101,
11'b11101110100,
11'b11101110101,
11'b11101110110,
11'b11110000101,
11'b11110000110: edge_mask_reg_512p7[432] <= 1'b1;
 		default: edge_mask_reg_512p7[432] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010111,
11'b110011000,
11'b110011001,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b10001000101,
11'b10001000110,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000100,
11'b10010000101,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000100,
11'b10110000101,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11010000101,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101,
11'b11101110100: edge_mask_reg_512p7[433] <= 1'b1;
 		default: edge_mask_reg_512p7[433] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110111,
11'b1010111000,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110100111,
11'b1110101000,
11'b10001000101,
11'b10001000110,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11010000100,
11'b11010000101,
11'b11010010100,
11'b11010010101,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101,
11'b11101110100,
11'b11101110101,
11'b11110000100: edge_mask_reg_512p7[434] <= 1'b1;
 		default: edge_mask_reg_512p7[434] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000111,
11'b10001000101,
11'b10001000110,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110101,
11'b10101110110,
11'b11001000100,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101: edge_mask_reg_512p7[435] <= 1'b1;
 		default: edge_mask_reg_512p7[435] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110011000,
11'b1110011001,
11'b10001000101,
11'b10001000110,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000101,
11'b10010000110,
11'b10101000101,
11'b10101000110,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000101,
11'b10110000110,
11'b11001000101,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101,
11'b11001110110,
11'b11010000101,
11'b11101010100,
11'b11101010101,
11'b11101100100,
11'b11101100101,
11'b11101110100,
11'b11101110101: edge_mask_reg_512p7[436] <= 1'b1;
 		default: edge_mask_reg_512p7[436] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1111101000,
11'b1111101001,
11'b10111110100,
11'b11011110100,
11'b11011110101: edge_mask_reg_512p7[437] <= 1'b1;
 		default: edge_mask_reg_512p7[437] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001001,
11'b110001010,
11'b110001011,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110101,
11'b1101110110,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001001,
11'b1110001010,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001110101,
11'b10001110110,
11'b10100110101,
11'b10100110110,
11'b10101000101,
11'b10101000110,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100101,
11'b10101100110,
11'b10101100111: edge_mask_reg_512p7[438] <= 1'b1;
 		default: edge_mask_reg_512p7[438] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111010,
11'b110111011,
11'b110111100,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010001101,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1100111010,
11'b1100111011,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b10001010110,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001011010,
11'b10001100110,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010011000,
11'b10010011001,
11'b10010011010,
11'b10010011011,
11'b10010101000,
11'b10101010110,
11'b10101010111,
11'b10101011000,
11'b10101100110,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110110,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b11001010111,
11'b11001011000,
11'b11001100110,
11'b11001100111,
11'b11001101000,
11'b11001110110,
11'b11001110111,
11'b11001111000,
11'b11010000110,
11'b11010000111,
11'b11010001000,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010100111,
11'b11101110110,
11'b11101110111,
11'b11110000110,
11'b11110000111,
11'b11110010111,
11'b11110011000: edge_mask_reg_512p7[439] <= 1'b1;
 		default: edge_mask_reg_512p7[439] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11001001,
11'b11001010,
11'b110111011,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1011001010,
11'b1011001011,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111001011,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111100110,
11'b10111100111,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b11011100110,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111110110: edge_mask_reg_512p7[440] <= 1'b1;
 		default: edge_mask_reg_512p7[440] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1101011010,
11'b1101011011,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10001111011,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10010001011,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10101101000,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110001001,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110011001,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110101001,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11010000110,
11'b11010000111,
11'b11010001000,
11'b11010001001,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010011001,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11101111000,
11'b11110000111,
11'b11110001000,
11'b11110010110,
11'b11110010111,
11'b11110011000: edge_mask_reg_512p7[441] <= 1'b1;
 		default: edge_mask_reg_512p7[441] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001001,
11'b111001010,
11'b111001011,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1101011001,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b10001100111,
11'b10001110110,
11'b10001110111,
11'b10001111000,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10101110101,
11'b10101110110,
11'b10101110111,
11'b10110000101,
11'b10110000110,
11'b10110000111,
11'b10110001000,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b11001110101,
11'b11001110110,
11'b11001110111,
11'b11010000101,
11'b11010000110,
11'b11010000111,
11'b11010010101,
11'b11010010110,
11'b11010010111,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110110,
11'b11010110111,
11'b11010111000: edge_mask_reg_512p7[442] <= 1'b1;
 		default: edge_mask_reg_512p7[442] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000111,
11'b10011001000,
11'b10011010111,
11'b10011011000,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b11010010110,
11'b11010010111,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000101,
11'b11011000110,
11'b11011000111,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11110110110,
11'b11111000101,
11'b11111000110,
11'b11111000111,
11'b11111010110: edge_mask_reg_512p7[443] <= 1'b1;
 		default: edge_mask_reg_512p7[443] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10110010110,
11'b10110010111,
11'b10110011000,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110101000,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b10110111000,
11'b10111000101,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b11010010110,
11'b11010010111,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110101,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000101,
11'b11011000110,
11'b11011000111,
11'b11110110101,
11'b11110110110,
11'b11111000101,
11'b11111000110: edge_mask_reg_512p7[444] <= 1'b1;
 		default: edge_mask_reg_512p7[444] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011100110,
11'b1011100111,
11'b1111100110,
11'b1111100111,
11'b10111110100,
11'b10111110101,
11'b11011110100: edge_mask_reg_512p7[445] <= 1'b1;
 		default: edge_mask_reg_512p7[445] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[446] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[447] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[448] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[449] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011010,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000101010,
11'b10000110111,
11'b10100000110,
11'b10100000111,
11'b10100001000,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100110110,
11'b10100110111,
11'b11000000110,
11'b11000000111,
11'b11000001000,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11000011000,
11'b11000100101,
11'b11000100110,
11'b11000100111,
11'b11100000110,
11'b11100000111,
11'b11100010110,
11'b11100100110: edge_mask_reg_512p7[450] <= 1'b1;
 		default: edge_mask_reg_512p7[450] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011001,
11'b1001011010,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011010,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000101010,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100110100,
11'b10100110101,
11'b10100110110,
11'b10100110111,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11000100100,
11'b11000100101,
11'b11000100110,
11'b11000100111,
11'b11000110101,
11'b11100100110: edge_mask_reg_512p7[451] <= 1'b1;
 		default: edge_mask_reg_512p7[451] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011010,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000101010,
11'b10000110111,
11'b10100000110,
11'b10100000111,
11'b10100001000,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100110110,
11'b10100110111,
11'b11000000101,
11'b11000000110,
11'b11000000111,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11000100101,
11'b11000100110,
11'b11000100111,
11'b11100000101,
11'b11100000110,
11'b11100010101,
11'b11100010110,
11'b11100100110: edge_mask_reg_512p7[452] <= 1'b1;
 		default: edge_mask_reg_512p7[452] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011010,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000101001,
11'b10000101010,
11'b10000110110,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10000111010,
11'b10000111011,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001001010,
11'b10001001011,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b10100101000,
11'b10100110110,
11'b10100110111,
11'b10100111000,
11'b10101000110,
11'b10101000111,
11'b10101001000,
11'b10101010111,
11'b10101011000,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11000100101,
11'b11000100110,
11'b11000100111,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010111,
11'b11001011000,
11'b11100100110,
11'b11100110110,
11'b11100110111,
11'b11101000110,
11'b11101000111: edge_mask_reg_512p7[453] <= 1'b1;
 		default: edge_mask_reg_512p7[453] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[454] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101010,
11'b10101011,
11'b100101010,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101011,
11'b110101100,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001011101,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001101101,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1100011010,
11'b1100011011,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b10000100111,
11'b10000101000,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10000111011,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001001011,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001011011,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101011,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111011,
11'b10100100111,
11'b10100101000,
11'b10100110111,
11'b10100111000,
11'b10100111001,
11'b10101000111,
11'b10101001000,
11'b10101001001,
11'b10101010111,
11'b10101011000,
11'b10101011001,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b10101111000,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010111,
11'b11001011000,
11'b11001100111,
11'b11001101000,
11'b11001110111,
11'b11001111000,
11'b11100110111,
11'b11101000110,
11'b11101000111,
11'b11101001000,
11'b11101010111,
11'b11101011000,
11'b11101100111,
11'b11101101000,
11'b11101110111,
11'b11101111000: edge_mask_reg_512p7[455] <= 1'b1;
 		default: edge_mask_reg_512p7[455] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101010,
11'b10101011,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001001101,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1100011010,
11'b1100011011,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110011010,
11'b10000100111,
11'b10000101000,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10000111011,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001001010,
11'b10001001011,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001011010,
11'b10001011011,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001101011,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10100100111,
11'b10100101000,
11'b10100110111,
11'b10100111000,
11'b10100111001,
11'b10101000111,
11'b10101001000,
11'b10101001001,
11'b10101010111,
11'b10101011000,
11'b10101100111,
11'b10101101000,
11'b10101110111,
11'b10101111000,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010111,
11'b11001011000,
11'b11001100111,
11'b11001101000,
11'b11001110111,
11'b11001111000,
11'b11100110110,
11'b11100110111,
11'b11101000110,
11'b11101000111,
11'b11101010111,
11'b11101100111,
11'b11101110111: edge_mask_reg_512p7[456] <= 1'b1;
 		default: edge_mask_reg_512p7[456] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[457] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111011,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010101010,
11'b1010101011,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101010,
11'b1110101011,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10001100111,
11'b10001101000,
11'b10001101001,
11'b10001101010,
11'b10001110111,
11'b10001111000,
11'b10001111001,
11'b10001111010,
11'b10010001000,
11'b10010001001,
11'b10010001010,
11'b10101010111,
11'b10101011000,
11'b10101011001,
11'b10101100111,
11'b10101101000,
11'b10101101001,
11'b10101110111,
11'b10101111000,
11'b10101111001,
11'b10101111010,
11'b10110001000,
11'b10110001001,
11'b10110001010,
11'b11001010111,
11'b11001011000,
11'b11001100111,
11'b11001101000,
11'b11001101001,
11'b11001110111,
11'b11001111000,
11'b11001111001,
11'b11010001000,
11'b11010001001,
11'b11101010111,
11'b11101011000,
11'b11101100111,
11'b11101101000,
11'b11101101001,
11'b11101110111,
11'b11101111000,
11'b11101111001,
11'b11110001000,
11'b11110001001: edge_mask_reg_512p7[458] <= 1'b1;
 		default: edge_mask_reg_512p7[458] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[459] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[460] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[461] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[462] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b100100110,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100100,
11'b1000100101,
11'b1000100110,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100100,
11'b1100100101,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b10000010100,
11'b10000010101,
11'b10000010110,
11'b10000100011,
11'b10000100100,
11'b10000100101,
11'b10000100110,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b10100100011,
11'b10100100100,
11'b10100100101,
11'b10100100110,
11'b11000010100,
11'b11000010101,
11'b11000100100,
11'b11000100101: edge_mask_reg_512p7[463] <= 1'b1;
 		default: edge_mask_reg_512p7[463] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b101000100,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010100,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b1000110100,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000011,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1100110011,
11'b1100110111,
11'b1100111000,
11'b1101000010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101010010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101000,
11'b1110101001,
11'b10001000011,
11'b10001000100,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100011,
11'b10010100100,
11'b10101100011,
11'b10101100100,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b10110000101,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100011,
11'b10110100100: edge_mask_reg_512p7[464] <= 1'b1;
 		default: edge_mask_reg_512p7[464] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100101,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100100,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b10001100011,
11'b10001100100,
11'b10001110011,
11'b10001110100,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10101110011,
11'b10110000011,
11'b10110000100,
11'b10110010011,
11'b10110010100: edge_mask_reg_512p7[465] <= 1'b1;
 		default: edge_mask_reg_512p7[465] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110011,
11'b1110110100,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b10001100011,
11'b10001100100,
11'b10001110011,
11'b10001110100,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100,
11'b10010110011,
11'b10101110011,
11'b10110000011,
11'b10110010011: edge_mask_reg_512p7[466] <= 1'b1;
 		default: edge_mask_reg_512p7[466] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000110,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1010110,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111001,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1101000111,
11'b1101001000,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110101000,
11'b10001010011,
11'b10001010100,
11'b10001100011,
11'b10001100100,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010011,
11'b10010010100,
11'b10101100011,
11'b10101100100,
11'b10101110011,
11'b10101110100,
11'b10110000011,
11'b10110000100: edge_mask_reg_512p7[467] <= 1'b1;
 		default: edge_mask_reg_512p7[467] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110100,
11'b1110110101,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011000,
11'b1111011001,
11'b10001100011,
11'b10001100100,
11'b10001110011,
11'b10001110100,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010110100,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10011000100,
11'b10011000101,
11'b10011000110,
11'b10101100011,
11'b10101110011,
11'b10101110100,
11'b10110000011,
11'b10110000100,
11'b10110010011,
11'b10110010100,
11'b10110010101,
11'b10110100011,
11'b10110100100,
11'b10110100101,
11'b10110110100,
11'b10110110101,
11'b10110110110,
11'b10111000101,
11'b11010010100,
11'b11010100100,
11'b11010100101,
11'b11010110100,
11'b11010110101: edge_mask_reg_512p7[468] <= 1'b1;
 		default: edge_mask_reg_512p7[468] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100110,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110110,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000110,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000111,
11'b111001000,
11'b111001001,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1011000111,
11'b1011001000,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110100010,
11'b1110100011,
11'b1110100100,
11'b1110100101,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110110010,
11'b1110110011,
11'b1110110100,
11'b1110110101,
11'b1110110111,
11'b1110111000,
11'b10001100011,
11'b10001100100,
11'b10001110011,
11'b10001110100,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010011,
11'b10010010100,
11'b10010100011,
11'b10010100100,
11'b10010110011,
11'b10010110100,
11'b10101110011,
11'b10110000011,
11'b10110010011: edge_mask_reg_512p7[469] <= 1'b1;
 		default: edge_mask_reg_512p7[469] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10111001,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000101,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101010101,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110100111,
11'b110101000,
11'b110101001,
11'b1000110100,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010011,
11'b1001010100,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1100110100,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110101000,
11'b10001000011,
11'b10001000100,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010010011,
11'b10010010100,
11'b10101000011,
11'b10101010011,
11'b10101010100,
11'b10101100011,
11'b10101100100,
11'b10101110011,
11'b10110000011: edge_mask_reg_512p7[470] <= 1'b1;
 		default: edge_mask_reg_512p7[470] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10110110,
11'b10110111,
11'b10111000,
11'b10111001,
11'b11000110,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110110110,
11'b110110111,
11'b110111000,
11'b110111001,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111010110,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010110110,
11'b1010110111,
11'b1010111000,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1111000100,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111001000,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111110111,
11'b1111111000,
11'b10011000011,
11'b10011000100,
11'b10011000101,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011010110,
11'b10011100100,
11'b10011100101,
11'b10011100110,
11'b10011110101,
11'b10011110110,
11'b10111000011,
11'b10111000100,
11'b10111000101,
11'b10111010011,
11'b10111010100,
11'b10111010101,
11'b10111100011,
11'b10111100100,
11'b10111100101,
11'b10111110100,
11'b10111110101,
11'b11011000100,
11'b11011010100,
11'b11011010101,
11'b11011100100,
11'b11011100101,
11'b11011110100,
11'b11011110101: edge_mask_reg_512p7[471] <= 1'b1;
 		default: edge_mask_reg_512p7[471] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010010111,
11'b10010011000,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011011000,
11'b10011011001,
11'b10110010111,
11'b10110011000,
11'b10110100111,
11'b10110101000,
11'b10110110111,
11'b10110111000,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b11010010111,
11'b11010011000,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11110010111,
11'b11110011000,
11'b11110100110,
11'b11110100111,
11'b11110101000,
11'b11110110110,
11'b11110110111,
11'b11110111000,
11'b11111000110,
11'b11111000111,
11'b11111001000,
11'b11111010110,
11'b11111010111,
11'b11111011000: edge_mask_reg_512p7[472] <= 1'b1;
 		default: edge_mask_reg_512p7[472] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1101111000,
11'b1101111001,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b10010000111,
11'b10010001000,
11'b10010001001,
11'b10010010111,
11'b10010011000,
11'b10010011001,
11'b10010100111,
11'b10010101000,
11'b10010101001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011011000,
11'b10011011001,
11'b10110000111,
11'b10110001000,
11'b10110010111,
11'b10110011000,
11'b10110100111,
11'b10110101000,
11'b10110110111,
11'b10110111000,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b11010000111,
11'b11010001000,
11'b11010010110,
11'b11010010111,
11'b11010011000,
11'b11010100110,
11'b11010100111,
11'b11010101000,
11'b11010110110,
11'b11010110111,
11'b11010111000,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11110000111,
11'b11110001000,
11'b11110010110,
11'b11110010111,
11'b11110011000,
11'b11110100110,
11'b11110100111,
11'b11110101000,
11'b11110110110,
11'b11110110111,
11'b11110111000,
11'b11111000110,
11'b11111000111,
11'b11111001000,
11'b11111010110,
11'b11111010111,
11'b11111011000: edge_mask_reg_512p7[473] <= 1'b1;
 		default: edge_mask_reg_512p7[473] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001010,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10110111,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11000111,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110110111,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b111000111,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111010111,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1011000111,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011010111,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1111000111,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111010110,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10010110111,
11'b10010111000,
11'b10010111001,
11'b10011000110,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011010110,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011100110,
11'b10011100111,
11'b10011101000,
11'b10011110110,
11'b10011110111,
11'b10110110111,
11'b10110111000,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010101,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100100,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110100,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b11010110111,
11'b11010111000,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010101,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100100,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011110100,
11'b11011110101,
11'b11011110110,
11'b11110110111,
11'b11110111000,
11'b11111000110,
11'b11111000111,
11'b11111001000,
11'b11111010101,
11'b11111010110,
11'b11111010111,
11'b11111011000,
11'b11111100101,
11'b11111100110,
11'b11111100111,
11'b11111110101,
11'b11111110110: edge_mask_reg_512p7[474] <= 1'b1;
 		default: edge_mask_reg_512p7[474] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[475] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[476] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000010111: edge_mask_reg_512p7[477] <= 1'b1;
 		default: edge_mask_reg_512p7[477] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011100111,
11'b1011101000: edge_mask_reg_512p7[478] <= 1'b1;
 		default: edge_mask_reg_512p7[478] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[479] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[480] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100111011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000101011,
11'b1000111011,
11'b1000111100,
11'b1001001100,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100101011,
11'b1100101100,
11'b1100111011,
11'b1100111100,
11'b10000010110,
11'b10000010111,
11'b10000011000: edge_mask_reg_512p7[481] <= 1'b1;
 		default: edge_mask_reg_512p7[481] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001010,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100111001,
11'b1100111010,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000100101,
11'b10000100110,
11'b10000100111,
11'b10100000110,
11'b10100010100,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100100110,
11'b11000000101,
11'b11000010101: edge_mask_reg_512p7[482] <= 1'b1;
 		default: edge_mask_reg_512p7[482] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1000011001,
11'b1000101001,
11'b1000101010,
11'b1100011001,
11'b1100011010,
11'b1100101001,
11'b1100101010,
11'b10000010110: edge_mask_reg_512p7[483] <= 1'b1;
 		default: edge_mask_reg_512p7[483] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001010,
11'b101001011,
11'b101001100,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1100010101,
11'b1100010110,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100110,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101001010,
11'b1101001011,
11'b10000010101,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011010,
11'b10000011011,
11'b10000100110,
11'b10000100111,
11'b10000101000,
11'b10000101010,
11'b10000101011,
11'b10100000110,
11'b10100000111,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100100101,
11'b10100100110,
11'b10100100111,
11'b11000000101,
11'b11000000110,
11'b11000010101,
11'b11000010110,
11'b11000100110: edge_mask_reg_512p7[484] <= 1'b1;
 		default: edge_mask_reg_512p7[484] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[485] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[486] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011100110,
11'b1011100111,
11'b1111100110,
11'b1111100111,
11'b10111110100,
11'b10111110101,
11'b11011110100: edge_mask_reg_512p7[487] <= 1'b1;
 		default: edge_mask_reg_512p7[487] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1011100110,
11'b1011100111,
11'b1111100110: edge_mask_reg_512p7[488] <= 1'b1;
 		default: edge_mask_reg_512p7[488] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10100110,
11'b10100111,
11'b10110101,
11'b10110110,
11'b10110111,
11'b10111000,
11'b11000110,
11'b11000111,
11'b11001000,
11'b110110101,
11'b110110110,
11'b110110111,
11'b110111000,
11'b111000101,
11'b111000110,
11'b111000111,
11'b111001000,
11'b111010101,
11'b111010110,
11'b111010111,
11'b111011000,
11'b1010110101,
11'b1010110110,
11'b1010110111,
11'b1011000101,
11'b1011000110,
11'b1011000111,
11'b1011010100,
11'b1011010101,
11'b1011010110,
11'b1011010111,
11'b1011011000,
11'b1011100101,
11'b1011100110,
11'b1011100111,
11'b1011101000,
11'b1111000101,
11'b1111000110,
11'b1111000111,
11'b1111010100,
11'b1111010101,
11'b1111010110,
11'b1111010111,
11'b1111100100,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111110111,
11'b10011000100,
11'b10011010011,
11'b10011010100,
11'b10011010101,
11'b10011100011,
11'b10011100100,
11'b10011100101,
11'b10111000011,
11'b10111000100,
11'b10111010011,
11'b10111010100,
11'b10111100011,
11'b10111100100,
11'b10111110100: edge_mask_reg_512p7[489] <= 1'b1;
 		default: edge_mask_reg_512p7[489] <= 1'b0;
 	endcase

    case({x,y,z})
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000111000,
11'b1000111001,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b10000011000,
11'b10000011001,
11'b10100001000,
11'b10100001001,
11'b10100011000,
11'b10100011001,
11'b11000001000,
11'b11000001001,
11'b11000011000,
11'b11000011001,
11'b11100001000,
11'b11100001001,
11'b11100011000,
11'b11100011001: edge_mask_reg_512p7[490] <= 1'b1;
 		default: edge_mask_reg_512p7[490] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111011,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1001010100,
11'b1001010101,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101010,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001111010,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010001010: edge_mask_reg_512p7[491] <= 1'b1;
 		default: edge_mask_reg_512p7[491] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001010,
11'b101001010,
11'b101001011,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b101111100,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001010,
11'b111001011,
11'b1001010100,
11'b1001010101,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1101111100,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110100100,
11'b1110100101,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001010,
11'b1111001011,
11'b10001110011,
11'b10001110100,
11'b10010000011,
11'b10010000100,
11'b10010000101,
11'b10010001010,
11'b10010001011,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010011010,
11'b10010011011,
11'b10010101011: edge_mask_reg_512p7[492] <= 1'b1;
 		default: edge_mask_reg_512p7[492] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10000110,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10010101,
11'b10010110,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10100101,
11'b10100110,
11'b10100111,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001010,
11'b101001010,
11'b101001011,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100100,
11'b101100101,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110011,
11'b101110100,
11'b101110101,
11'b101110110,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110000011,
11'b110000100,
11'b110000101,
11'b110000110,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110010011,
11'b110010100,
11'b110010101,
11'b110010110,
11'b110010111,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110100011,
11'b110100100,
11'b110100101,
11'b110100110,
11'b110100111,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110110100,
11'b110110101,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b1001010100,
11'b1001010101,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100011,
11'b1001100100,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110010,
11'b1001110011,
11'b1001110100,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000010,
11'b1010000011,
11'b1010000100,
11'b1010000101,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010011,
11'b1010010100,
11'b1010010101,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010100011,
11'b1010100100,
11'b1010100101,
11'b1010100110,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010110011,
11'b1010110100,
11'b1010110101,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100010,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110010,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000010,
11'b1110000011,
11'b1110000100,
11'b1110000101,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010010,
11'b1110010011,
11'b1110010100,
11'b1110010101,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100010,
11'b1110100100,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111001,
11'b1110111010,
11'b10001110011: edge_mask_reg_512p7[493] <= 1'b1;
 		default: edge_mask_reg_512p7[493] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111001,
11'b100101001,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001011,
11'b1000010111,
11'b1000011000,
11'b1000011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1100010111,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b10000010110,
11'b10000010111,
11'b10000011000,
11'b10000011010,
11'b10000100111,
11'b10000101000,
11'b10100000110,
11'b10100000111,
11'b10100001000,
11'b10100010101,
11'b10100010110,
11'b10100010111,
11'b10100011000,
11'b10100100111,
11'b11000000101,
11'b11000000110,
11'b11000000111,
11'b11000010101,
11'b11000010110,
11'b11000010111,
11'b11100000110,
11'b11100010110: edge_mask_reg_512p7[494] <= 1'b1;
 		default: edge_mask_reg_512p7[494] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[495] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[496] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[497] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001001,
11'b1001010,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111001,
11'b1111010,
11'b1111011,
11'b100101010,
11'b100111001,
11'b100111010,
11'b100111011,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101001100,
11'b101011010,
11'b101011011,
11'b101011100,
11'b101101010,
11'b101101011,
11'b101101100,
11'b101111010,
11'b101111011,
11'b101111100,
11'b1000011001,
11'b1000101001,
11'b1000101010,
11'b1000101011,
11'b1000111001,
11'b1000111010,
11'b1000111011,
11'b1000111100,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001001100,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001011100,
11'b1001101010,
11'b1001101011,
11'b1001101100,
11'b1001111010,
11'b1001111011,
11'b1001111100,
11'b1100011000,
11'b1100011001,
11'b1100011010,
11'b1100011011,
11'b1100101000,
11'b1100101001,
11'b1100101010,
11'b1100101011,
11'b1100101100,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1100111011,
11'b1100111100,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101001011,
11'b1101001100,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101011100,
11'b1101101010,
11'b1101101011,
11'b1101101100,
11'b10000010111,
11'b10000011000,
11'b10000011001,
11'b10000011011,
11'b10000100111,
11'b10000101000,
11'b10000101001,
11'b10000101011,
11'b10000110111,
11'b10000111000,
11'b10000111001,
11'b10000111011,
11'b10001000111,
11'b10001001000,
11'b10001001001,
11'b10001001011,
11'b10001010111,
11'b10001011000,
11'b10001011001,
11'b10100010111,
11'b10100011000,
11'b10100100111,
11'b10100101000,
11'b10100101001,
11'b10100110111,
11'b10100111000,
11'b10100111001,
11'b10101000111,
11'b10101001000,
11'b10101001001,
11'b10101010111,
11'b10101011000,
11'b11000010111,
11'b11000011000,
11'b11000100110,
11'b11000100111,
11'b11000101000,
11'b11000110110,
11'b11000110111,
11'b11000111000,
11'b11001000110,
11'b11001000111,
11'b11001001000,
11'b11001010111,
11'b11001011000,
11'b11100010111,
11'b11100100110,
11'b11100100111,
11'b11100110111,
11'b11101000111: edge_mask_reg_512p7[498] <= 1'b1;
 		default: edge_mask_reg_512p7[498] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1111010,
11'b1111011,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001001,
11'b11001010,
11'b101111011,
11'b101111100,
11'b110001010,
11'b110001011,
11'b110001100,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1010001010,
11'b1010001011,
11'b1010001100,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010011101,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010101101,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101001,
11'b1011101010,
11'b1110001010,
11'b1110001011,
11'b1110001100,
11'b1110011010,
11'b1110011011,
11'b1110011100,
11'b1110101010,
11'b1110101011,
11'b1110101100,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1110111100,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b10010101001,
11'b10010101010,
11'b10010101011,
11'b10010111001,
11'b10010111010,
11'b10010111011,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011011001,
11'b10011011010,
11'b10011101001,
11'b10011101010,
11'b10110101001,
11'b10110101010,
11'b10110111001,
11'b10110111010,
11'b10111001001,
11'b10111001010,
11'b10111011001,
11'b10111011010,
11'b10111101000,
11'b10111101001,
11'b10111101010,
11'b11010101001,
11'b11010101010,
11'b11010111001,
11'b11010111010,
11'b11011001000,
11'b11011001001,
11'b11011001010,
11'b11011011000,
11'b11011011001,
11'b11011011010,
11'b11011101000,
11'b11011101001,
11'b11110101000,
11'b11110101001,
11'b11110101010,
11'b11110111000,
11'b11110111001,
11'b11110111010,
11'b11111001000,
11'b11111001001,
11'b11111001010,
11'b11111011000,
11'b11111011001,
11'b11111101000,
11'b11111101001: edge_mask_reg_512p7[499] <= 1'b1;
 		default: edge_mask_reg_512p7[499] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110101010,
11'b1110101011,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111001100,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111011100,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10011101010,
11'b10011101011,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111101001,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b11011000111,
11'b11011001000,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011101000,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111010110,
11'b11111010111,
11'b11111100101,
11'b11111100110,
11'b11111100111: edge_mask_reg_512p7[500] <= 1'b1;
 		default: edge_mask_reg_512p7[500] <= 1'b0;
 	endcase

    case({x,y,z})
11'b10001010,
11'b10001011,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001000,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1010011010,
11'b1010011011,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001000,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011001100,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1011011100,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001000,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111010111,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111011011,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111101011,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10010111000,
11'b10010111001,
11'b10011000111,
11'b10011001000,
11'b10011001001,
11'b10011001010,
11'b10011001011,
11'b10011010111,
11'b10011011000,
11'b10011011001,
11'b10011011010,
11'b10011011011,
11'b10011100111,
11'b10011101000,
11'b10011101001,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10110110111,
11'b10110111000,
11'b10110111001,
11'b10111000110,
11'b10111000111,
11'b10111001000,
11'b10111001001,
11'b10111010110,
11'b10111010111,
11'b10111011000,
11'b10111011001,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111101000,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b10111111000,
11'b11010110111,
11'b11010111000,
11'b11011000110,
11'b11011000111,
11'b11011001000,
11'b11011010110,
11'b11011010111,
11'b11011011000,
11'b11011100101,
11'b11011100110,
11'b11011100111,
11'b11011101000,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111000110,
11'b11111000111,
11'b11111010110,
11'b11111010111,
11'b11111100101,
11'b11111100110: edge_mask_reg_512p7[501] <= 1'b1;
 		default: edge_mask_reg_512p7[501] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[502] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[503] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[504] <= 1'b0;
 	endcase

    case({x,y,z})
11'b101001100,
11'b101011100,
11'b101101100,
11'b101111100,
11'b110001100,
11'b110011100,
11'b110101100,
11'b110111100,
11'b1001001100,
11'b1001001101,
11'b1001011100,
11'b1001011101,
11'b1001101100,
11'b1001101101,
11'b1001111100,
11'b1001111101,
11'b1010001100,
11'b1010001101,
11'b1010011100,
11'b1010011101,
11'b1010101100,
11'b1010101101,
11'b1010111100,
11'b1010111101,
11'b1011001100,
11'b1101001100,
11'b1101001101,
11'b1101011100,
11'b1101011101,
11'b1101101100,
11'b1101101101,
11'b1101111011,
11'b1101111100,
11'b1101111101,
11'b1110001011,
11'b1110001100,
11'b1110001101,
11'b1110011011,
11'b1110011100,
11'b1110011101,
11'b1110101100,
11'b1110101101,
11'b1110111100,
11'b1110111101,
11'b1111001100,
11'b1111001101,
11'b10001101011,
11'b10001111011,
11'b10001111100,
11'b10001111101,
11'b10001111110,
11'b10010001010,
11'b10010001011,
11'b10010001100,
11'b10010001101,
11'b10010001110,
11'b10010011010,
11'b10010011011,
11'b10010011100,
11'b10010011101,
11'b10010011110,
11'b10010101011,
11'b10010101100,
11'b10010101101,
11'b10010111100,
11'b10010111101,
11'b10011001100,
11'b10011001101,
11'b10101101011,
11'b10101111010,
11'b10101111011,
11'b10101111100,
11'b10110001010,
11'b10110001011,
11'b10110001100,
11'b10110001101,
11'b10110011010,
11'b10110011011,
11'b10110011100,
11'b10110011101,
11'b10110101011,
11'b10110101100,
11'b10110101101,
11'b10110111011,
11'b10110111100,
11'b10110111101,
11'b10111001100,
11'b10111001101,
11'b11001111010,
11'b11001111011,
11'b11001111100,
11'b11010001010,
11'b11010001011,
11'b11010001100,
11'b11010011010,
11'b11010011011,
11'b11010011100,
11'b11010011101,
11'b11010101011,
11'b11010101100,
11'b11010101101,
11'b11010111011,
11'b11010111100,
11'b11101111001,
11'b11101111010,
11'b11101111011,
11'b11110001010,
11'b11110001011,
11'b11110001100,
11'b11110011010,
11'b11110011011,
11'b11110011100,
11'b11110101011,
11'b11110101100,
11'b11110111011,
11'b11110111100: edge_mask_reg_512p7[505] <= 1'b1;
 		default: edge_mask_reg_512p7[505] <= 1'b0;
 	endcase

    case({x,y,z})
11'b110111,
11'b111000,
11'b111001,
11'b1000111,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10000111,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10010111,
11'b10011000,
11'b10011001,
11'b10011010,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b110000111,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110011001,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1100101001,
11'b1100110110,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1110001000,
11'b1110001001,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10010000011,
11'b10010000100,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10110000011,
11'b10110000100,
11'b11001000101,
11'b11001000110,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101,
11'b11001100110,
11'b11001110100,
11'b11001110101: edge_mask_reg_512p7[506] <= 1'b1;
 		default: edge_mask_reg_512p7[506] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001001,
11'b1001010,
11'b1010111,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1100111,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1110111,
11'b1111000,
11'b1111001,
11'b1111010,
11'b10001001,
11'b10001010,
11'b100100111,
11'b100101000,
11'b100101001,
11'b100101010,
11'b100110110,
11'b100110111,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101000110,
11'b101000111,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101111000,
11'b101111001,
11'b101111010,
11'b1000100101,
11'b1000100111,
11'b1000101000,
11'b1000101001,
11'b1000101010,
11'b1000110100,
11'b1000110101,
11'b1000110110,
11'b1000110111,
11'b1000111000,
11'b1000111001,
11'b1000111010,
11'b1001000100,
11'b1001000101,
11'b1001000110,
11'b1001000111,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001001011,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1100100100,
11'b1100100101,
11'b1100100111,
11'b1100101000,
11'b1100101001,
11'b1100110011,
11'b1100110100,
11'b1100110101,
11'b1100110110,
11'b1100110111,
11'b1100111000,
11'b1100111001,
11'b1100111010,
11'b1101000011,
11'b1101000100,
11'b1101000101,
11'b1101000110,
11'b1101000111,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010011,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101100011,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101111001,
11'b10000110011,
11'b10000110100,
11'b10000110101,
11'b10000110110,
11'b10001000011,
11'b10001000100,
11'b10001000101,
11'b10001000110,
11'b10001000111,
11'b10001010011,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001010111,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10100110100,
11'b10100110101,
11'b10101000011,
11'b10101000100,
11'b10101000101,
11'b10101000110,
11'b10101000111,
11'b10101010011,
11'b10101010100,
11'b10101010101,
11'b10101010110,
11'b10101010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b11001000101,
11'b11001000110,
11'b11001010100,
11'b11001010101,
11'b11001010110,
11'b11001100100,
11'b11001100101: edge_mask_reg_512p7[507] <= 1'b1;
 		default: edge_mask_reg_512p7[507] <= 1'b0;
 	endcase

    case({x,y,z})
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b11001000,
11'b11001001,
11'b11001010,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110011100,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b110101100,
11'b110111000,
11'b110111001,
11'b110111010,
11'b110111011,
11'b110111100,
11'b111001001,
11'b111001010,
11'b111001011,
11'b111011001,
11'b111011010,
11'b1001011001,
11'b1001011010,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010110,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010011100,
11'b1010100111,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1010101100,
11'b1010110111,
11'b1010111000,
11'b1010111001,
11'b1010111010,
11'b1010111011,
11'b1010111100,
11'b1011001001,
11'b1011001010,
11'b1011001011,
11'b1011011001,
11'b1011011010,
11'b1011011011,
11'b1101100110,
11'b1101101001,
11'b1101101010,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010101,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110100110,
11'b1110100111,
11'b1110101000,
11'b1110101001,
11'b1110101010,
11'b1110101011,
11'b1110110110,
11'b1110110111,
11'b1110111000,
11'b1110111001,
11'b1110111010,
11'b1110111011,
11'b1111001001,
11'b1111001010,
11'b1111001011,
11'b1111011001,
11'b1111011010,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010001000,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10010011000,
11'b10010100100,
11'b10010100101,
11'b10010100110,
11'b10010100111,
11'b10010101000,
11'b10010110101,
11'b10010110110,
11'b10010110111,
11'b10010111000,
11'b10101110101,
11'b10101110110,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110,
11'b10110010111,
11'b10110100100,
11'b10110100101,
11'b10110100110,
11'b10110100111,
11'b10110110101,
11'b10110110110,
11'b10110110111,
11'b11010000100,
11'b11010000101,
11'b11010010101,
11'b11010010110,
11'b11010100101,
11'b11010100110,
11'b11010100111,
11'b11010110101,
11'b11010110110,
11'b11010110111: edge_mask_reg_512p7[508] <= 1'b1;
 		default: edge_mask_reg_512p7[508] <= 1'b0;
 	endcase

    case({x,y,z})
11'b111000,
11'b111001,
11'b1001000,
11'b1001001,
11'b1001010,
11'b1011000,
11'b1011001,
11'b1011010,
11'b1011011,
11'b1101000,
11'b1101001,
11'b1101010,
11'b1101011,
11'b1111000,
11'b1111001,
11'b1111010,
11'b1111011,
11'b10001000,
11'b10001001,
11'b10001010,
11'b10001011,
11'b10011000,
11'b10011001,
11'b10011010,
11'b10011011,
11'b10101000,
11'b10101001,
11'b10101010,
11'b10101011,
11'b10111000,
11'b10111001,
11'b10111010,
11'b10111011,
11'b100111000,
11'b100111001,
11'b100111010,
11'b101001000,
11'b101001001,
11'b101001010,
11'b101001011,
11'b101010110,
11'b101010111,
11'b101011000,
11'b101011001,
11'b101011010,
11'b101011011,
11'b101100110,
11'b101100111,
11'b101101000,
11'b101101001,
11'b101101010,
11'b101101011,
11'b101110111,
11'b101111000,
11'b101111001,
11'b101111010,
11'b101111011,
11'b110001000,
11'b110001001,
11'b110001010,
11'b110001011,
11'b110011000,
11'b110011001,
11'b110011010,
11'b110011011,
11'b110101000,
11'b110101001,
11'b110101010,
11'b110101011,
11'b1000111010,
11'b1001001000,
11'b1001001001,
11'b1001001010,
11'b1001010101,
11'b1001010110,
11'b1001010111,
11'b1001011000,
11'b1001011001,
11'b1001011010,
11'b1001011011,
11'b1001100101,
11'b1001100110,
11'b1001100111,
11'b1001101000,
11'b1001101001,
11'b1001101010,
11'b1001101011,
11'b1001110101,
11'b1001110110,
11'b1001110111,
11'b1001111000,
11'b1001111001,
11'b1001111010,
11'b1001111011,
11'b1010000110,
11'b1010000111,
11'b1010001000,
11'b1010001001,
11'b1010001010,
11'b1010001011,
11'b1010010111,
11'b1010011000,
11'b1010011001,
11'b1010011010,
11'b1010011011,
11'b1010101000,
11'b1010101001,
11'b1010101010,
11'b1010101011,
11'b1101000101,
11'b1101001000,
11'b1101001001,
11'b1101001010,
11'b1101010100,
11'b1101010101,
11'b1101010110,
11'b1101010111,
11'b1101011000,
11'b1101011001,
11'b1101011010,
11'b1101011011,
11'b1101100011,
11'b1101100100,
11'b1101100101,
11'b1101100110,
11'b1101100111,
11'b1101101000,
11'b1101101001,
11'b1101101010,
11'b1101101011,
11'b1101110011,
11'b1101110100,
11'b1101110101,
11'b1101110110,
11'b1101110111,
11'b1101111000,
11'b1101111001,
11'b1101111010,
11'b1101111011,
11'b1110000100,
11'b1110000101,
11'b1110000110,
11'b1110000111,
11'b1110001000,
11'b1110001001,
11'b1110001010,
11'b1110001011,
11'b1110010110,
11'b1110010111,
11'b1110011000,
11'b1110011001,
11'b1110011010,
11'b1110011011,
11'b1110101001,
11'b1110101010,
11'b10001000101,
11'b10001010100,
11'b10001010101,
11'b10001010110,
11'b10001100011,
11'b10001100100,
11'b10001100101,
11'b10001100110,
11'b10001100111,
11'b10001110011,
11'b10001110100,
11'b10001110101,
11'b10001110110,
11'b10001110111,
11'b10010000100,
11'b10010000101,
11'b10010000110,
11'b10010000111,
11'b10010010100,
11'b10010010101,
11'b10010010110,
11'b10010010111,
11'b10101100011,
11'b10101100100,
11'b10101100101,
11'b10101100110,
11'b10101110011,
11'b10101110100,
11'b10101110101,
11'b10101110110,
11'b10110000100,
11'b10110000101,
11'b10110000110,
11'b10110010100,
11'b10110010101,
11'b10110010110: edge_mask_reg_512p7[509] <= 1'b1;
 		default: edge_mask_reg_512p7[509] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p7[510] <= 1'b0;
 	endcase

    case({x,y,z})
11'b11001000,
11'b111001001,
11'b111001010,
11'b111011000,
11'b111011001,
11'b111011010,
11'b1011011000,
11'b1011011001,
11'b1011011010,
11'b1011100111,
11'b1011101000,
11'b1011101001,
11'b1011101010,
11'b1111011000,
11'b1111011001,
11'b1111011010,
11'b1111100101,
11'b1111100110,
11'b1111100111,
11'b1111101000,
11'b1111101001,
11'b1111101010,
11'b1111110111,
11'b1111111000,
11'b1111111001,
11'b10011100101,
11'b10011100110,
11'b10011100111,
11'b10011110101,
11'b10011110110,
11'b10011110111,
11'b10011111000,
11'b10111100101,
11'b10111100110,
11'b10111100111,
11'b10111110101,
11'b10111110110,
11'b10111110111,
11'b11011100101,
11'b11011100110,
11'b11011110100,
11'b11011110101,
11'b11011110110,
11'b11011110111,
11'b11111110101,
11'b11111110110: edge_mask_reg_512p7[511] <= 1'b1;
 		default: edge_mask_reg_512p7[511] <= 1'b0;
 	endcase

end
endmodule

