/*******************************************
****** Wuhan university of technology ******
****** Ruige Lee ******
year: 2019
month: 3
date: 4
hour: 17
minutes: 3
second: 59
********************************************/

module prm_LUTX1_Po_4_5_4_chk512p3(
	input [3:0] x,
	input [4:0] y,
	input [3:0] z,
	output [511:0] edge_mask_512p3
);

	reg [511:0] edge_mask_reg_512p3;
	assign edge_mask_512p3= edge_mask_reg_512p3;

always @( *) begin
    case({x,y,z})
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010000,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110000,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110000,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100110111,
13'b101100111000,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101101000,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101111000,
13'b111101111001,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000111,
13'b111111001000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010111,
13'b111111011000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100111,
13'b111111101000,
13'b1000101010010,
13'b1000101010011,
13'b1000101100010,
13'b1000101100011,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100010,
13'b1000110100011,
13'b1000110110010,
13'b1000110110011: edge_mask_reg_512p3[0] <= 1'b1;
 		default: edge_mask_reg_512p3[0] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101111000,
13'b100101111001,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101111000,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110001000,
13'b110110001001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110111000,
13'b111110111001,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100111,
13'b111111101000,
13'b1000110010011,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1001111000011,
13'b1001111010011: edge_mask_reg_512p3[1] <= 1'b1;
 		default: edge_mask_reg_512p3[1] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100010110,
13'b1100010111,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11100100110,
13'b11100100111,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110000,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000000,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110000,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100100111,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000001,
13'b101101000010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110100110110,
13'b110100110111,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101000001,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100110,
13'b111101100111,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100111,
13'b111110101000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110111,
13'b111110111000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000111,
13'b111111001000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010111,
13'b111111011000,
13'b111111100001,
13'b111111100010,
13'b111111100111,
13'b111111101000,
13'b1000101100001,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110010001,
13'b1000110010010,
13'b1000110100001,
13'b1000110100010,
13'b1000110110001,
13'b1000110110010: edge_mask_reg_512p3[2] <= 1'b1;
 		default: edge_mask_reg_512p3[2] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100110000111,
13'b100110001000,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101110000111,
13'b101110001000,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110010111,
13'b110110011000,
13'b110110100010,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000111,
13'b111111001000,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000111010011,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100: edge_mask_reg_512p3[3] <= 1'b1;
 		default: edge_mask_reg_512p3[3] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101101000,
13'b10101101001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101111000,
13'b101101111001,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110001000,
13'b110110001001,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100111,
13'b111111101000,
13'b1000110010011,
13'b1000110010100,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1001110100011,
13'b1001110100100,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111100001,
13'b1001111100011,
13'b1010111000100,
13'b1010111010100: edge_mask_reg_512p3[4] <= 1'b1;
 		default: edge_mask_reg_512p3[4] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100100111001,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011001,
13'b101111011010,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b111101111000,
13'b111101111001,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b1000101111000,
13'b1000101111001,
13'b1000101111010,
13'b1000110001000,
13'b1000110001001,
13'b1000110001010,
13'b1000110001011,
13'b1000110011000,
13'b1000110011001,
13'b1000110011010,
13'b1000110011011,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110101010,
13'b1000110111000,
13'b1000110111001,
13'b1000110111010,
13'b1001101111000,
13'b1001101111001,
13'b1001101111010,
13'b1001110001000,
13'b1001110001001,
13'b1001110001010,
13'b1001110001011,
13'b1001110010111,
13'b1001110011000,
13'b1001110011001,
13'b1001110011010,
13'b1001110011011,
13'b1001110100111,
13'b1001110101000,
13'b1001110101001,
13'b1001110101010,
13'b1001110111000,
13'b1001110111001,
13'b1001110111010,
13'b1010101110111,
13'b1010101111000,
13'b1010101111001,
13'b1010101111010,
13'b1010110000111,
13'b1010110001000,
13'b1010110001001,
13'b1010110001010,
13'b1010110001011,
13'b1010110010111,
13'b1010110011000,
13'b1010110011001,
13'b1010110011010,
13'b1010110011011,
13'b1010110100111,
13'b1010110101000,
13'b1010110101001,
13'b1010110101010,
13'b1010110111000,
13'b1010110111001,
13'b1010110111010,
13'b1011101110111,
13'b1011101111000,
13'b1011101111001,
13'b1011110000111,
13'b1011110001000,
13'b1011110001001,
13'b1011110001010,
13'b1011110001011,
13'b1011110010111,
13'b1011110011000,
13'b1011110011001,
13'b1011110011010,
13'b1011110011011,
13'b1011110100111,
13'b1011110101000,
13'b1011110101001,
13'b1011110101010,
13'b1011110111000,
13'b1011110111001,
13'b1011110111010,
13'b1100101110111,
13'b1100101111000,
13'b1100101111001,
13'b1100110000111,
13'b1100110001000,
13'b1100110001001,
13'b1100110001010,
13'b1100110010111,
13'b1100110011000,
13'b1100110011001,
13'b1100110011010,
13'b1100110011011,
13'b1100110100111,
13'b1100110101000,
13'b1100110101001,
13'b1100110101010,
13'b1100110101011,
13'b1100110111000,
13'b1100110111001,
13'b1100110111010,
13'b1101101110111,
13'b1101101111000,
13'b1101101111001,
13'b1101110000111,
13'b1101110001000,
13'b1101110001001,
13'b1101110001010,
13'b1101110010111,
13'b1101110011000,
13'b1101110011001,
13'b1101110011010,
13'b1101110011011,
13'b1101110100111,
13'b1101110101000,
13'b1101110101001,
13'b1101110101010,
13'b1101110101011,
13'b1101110111000,
13'b1101110111001,
13'b1101110111010,
13'b1110101110111,
13'b1110101111000,
13'b1110101111001,
13'b1110110000111,
13'b1110110001000,
13'b1110110001001,
13'b1110110001010,
13'b1110110010110,
13'b1110110010111,
13'b1110110011000,
13'b1110110011001,
13'b1110110011010,
13'b1110110100111,
13'b1110110101000,
13'b1110110101001,
13'b1110110101010,
13'b1110110111000,
13'b1110110111001,
13'b1111110000110,
13'b1111110000111,
13'b1111110001000,
13'b1111110001001,
13'b1111110010110,
13'b1111110010111,
13'b1111110011000,
13'b1111110011001,
13'b1111110011010,
13'b1111110100111,
13'b1111110101000,
13'b1111110101001,
13'b1111110101010: edge_mask_reg_512p3[5] <= 1'b1;
 		default: edge_mask_reg_512p3[5] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10011111010,
13'b10011111011,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11011111010,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101100111010,
13'b101100111011,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001001,
13'b101111001010,
13'b101111011010,
13'b110101001010,
13'b110101001011,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b111100111010,
13'b111100111011,
13'b111101001010,
13'b111101001011,
13'b111101011010,
13'b111101011011,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110111001,
13'b111110111010,
13'b1000100111010,
13'b1000100111011,
13'b1000101001010,
13'b1000101001011,
13'b1000101011010,
13'b1000101011011,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1000110001001,
13'b1000110001010,
13'b1000110001011,
13'b1000110011001,
13'b1000110011010,
13'b1000110011011,
13'b1000110101001,
13'b1000110101010,
13'b1000110101011,
13'b1000110111001,
13'b1000110111010,
13'b1001100111010,
13'b1001100111011,
13'b1001101001010,
13'b1001101001011,
13'b1001101011010,
13'b1001101011011,
13'b1001101101001,
13'b1001101101010,
13'b1001101101011,
13'b1001101111001,
13'b1001101111010,
13'b1001101111011,
13'b1001110001001,
13'b1001110001010,
13'b1001110001011,
13'b1001110011001,
13'b1001110011010,
13'b1001110011011,
13'b1001110101001,
13'b1001110101010,
13'b1001110101011,
13'b1001110111001,
13'b1001110111010,
13'b1010100111010,
13'b1010100111011,
13'b1010101001010,
13'b1010101001011,
13'b1010101001100,
13'b1010101011010,
13'b1010101011011,
13'b1010101011100,
13'b1010101101001,
13'b1010101101010,
13'b1010101101011,
13'b1010101101100,
13'b1010101111001,
13'b1010101111010,
13'b1010101111011,
13'b1010110001001,
13'b1010110001010,
13'b1010110001011,
13'b1010110011001,
13'b1010110011010,
13'b1010110011011,
13'b1010110101001,
13'b1010110101010,
13'b1010110101011,
13'b1010110111001,
13'b1010110111010,
13'b1011100111010,
13'b1011100111011,
13'b1011100111100,
13'b1011101001010,
13'b1011101001011,
13'b1011101001100,
13'b1011101011010,
13'b1011101011011,
13'b1011101011100,
13'b1011101101001,
13'b1011101101010,
13'b1011101101011,
13'b1011101101100,
13'b1011101111001,
13'b1011101111010,
13'b1011101111011,
13'b1011101111100,
13'b1011110001001,
13'b1011110001010,
13'b1011110001011,
13'b1011110011001,
13'b1011110011010,
13'b1011110011011,
13'b1011110101001,
13'b1011110101010,
13'b1011110101011,
13'b1011110111001,
13'b1011110111010,
13'b1100100111010,
13'b1100100111011,
13'b1100101001010,
13'b1100101001011,
13'b1100101001100,
13'b1100101011010,
13'b1100101011011,
13'b1100101011100,
13'b1100101101001,
13'b1100101101010,
13'b1100101101011,
13'b1100101101100,
13'b1100101111001,
13'b1100101111010,
13'b1100101111011,
13'b1100101111100,
13'b1100110001001,
13'b1100110001010,
13'b1100110001011,
13'b1100110011001,
13'b1100110011010,
13'b1100110011011,
13'b1100110101001,
13'b1100110101010,
13'b1100110101011,
13'b1100110111001,
13'b1100110111010,
13'b1101101001010,
13'b1101101001011,
13'b1101101001100,
13'b1101101011010,
13'b1101101011011,
13'b1101101011100,
13'b1101101101001,
13'b1101101101010,
13'b1101101101011,
13'b1101101101100,
13'b1101101111001,
13'b1101101111010,
13'b1101101111011,
13'b1101110001001,
13'b1101110001010,
13'b1101110001011,
13'b1101110011001,
13'b1101110011010,
13'b1101110011011,
13'b1101110101001,
13'b1101110101010,
13'b1101110101011,
13'b1101110111001,
13'b1101110111010,
13'b1110101001010,
13'b1110101001011,
13'b1110101011010,
13'b1110101011011,
13'b1110101011100,
13'b1110101101010,
13'b1110101101011,
13'b1110101101100,
13'b1110101111001,
13'b1110101111010,
13'b1110101111011,
13'b1110110001001,
13'b1110110001010,
13'b1110110001011,
13'b1110110011001,
13'b1110110011010,
13'b1110110011011,
13'b1110110101001,
13'b1110110101010,
13'b1111101001011,
13'b1111101011010,
13'b1111101011011,
13'b1111101011100,
13'b1111101101010,
13'b1111101101011,
13'b1111101101100,
13'b1111101111001,
13'b1111101111010,
13'b1111101111011,
13'b1111110001001,
13'b1111110001010,
13'b1111110001011,
13'b1111110011001,
13'b1111110011010,
13'b1111110101000,
13'b1111110101001,
13'b1111110101010: edge_mask_reg_512p3[6] <= 1'b1;
 		default: edge_mask_reg_512p3[6] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100010110,
13'b1100010111,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100100100110,
13'b100100100111,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101100100111,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000010,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100110,
13'b111110100111,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110110,
13'b111110110111,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000110,
13'b111111000111,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010110,
13'b111111010111,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100110,
13'b111111100111,
13'b1000101010001,
13'b1000101010010,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1001101100001,
13'b1001101100010,
13'b1001101110001,
13'b1001101110010,
13'b1001110000001,
13'b1001110000010,
13'b1001110010001,
13'b1001110010010,
13'b1001110100001,
13'b1001110100010,
13'b1001110110001,
13'b1001111000001,
13'b1001111010001: edge_mask_reg_512p3[7] <= 1'b1;
 		default: edge_mask_reg_512p3[7] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100100100110,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101100100110,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111101000010,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010110,
13'b111110010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100110,
13'b111110100111,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110110,
13'b111110110111,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000110,
13'b111111000111,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010110,
13'b111111010111,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100110,
13'b111111100111,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1001101010000,
13'b1001101010001,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001111000000,
13'b1001111000001,
13'b1001111010000,
13'b1001111010001,
13'b1001111100000,
13'b1001111100001,
13'b1010101110000,
13'b1010101110001,
13'b1010110000001,
13'b1010110010001: edge_mask_reg_512p3[8] <= 1'b1;
 		default: edge_mask_reg_512p3[8] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000000,
13'b11110000001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110000,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100101,
13'b111110100110,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100110,
13'b111111100111,
13'b1000110110000,
13'b1000110110001,
13'b1000111000000,
13'b1000111000001,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010: edge_mask_reg_512p3[9] <= 1'b1;
 		default: edge_mask_reg_512p3[9] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[10] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010010,
13'b10010011,
13'b10010100,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100010,
13'b10100011,
13'b10100100,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110010,
13'b10110011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000010,
13'b11000011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11111001,
13'b1001100010,
13'b1001100011,
13'b1001100100,
13'b1001100101,
13'b1001100110,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001110010,
13'b1001110011,
13'b1001110100,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010000010,
13'b1010000011,
13'b1010000100,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010010001,
13'b1010010010,
13'b1010010011,
13'b1010010100,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010100001,
13'b1010100010,
13'b1010100011,
13'b1010100100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010110010,
13'b1010110011,
13'b1010110100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000010,
13'b1011000011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b10001010011,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100010,
13'b10001100011,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001110010,
13'b10001110011,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010000010,
13'b10010000011,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010010001,
13'b10010010010,
13'b10010010011,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010100010,
13'b10010100011,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010110010,
13'b10010110011,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000010,
13'b10011000011,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101001,
13'b10011101010,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110010,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010000010,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b100000111001,
13'b100000111010,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000011,
13'b100011000100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b101001001001,
13'b101001001010,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001011001,
13'b101001011010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111001,
13'b101010111010,
13'b101011001001,
13'b101011001010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110100,
13'b111010110101,
13'b1000001110100,
13'b1000001110101,
13'b1000010000100,
13'b1000010000101,
13'b1000010010100,
13'b1000010010101,
13'b1000010100100,
13'b1000010100101: edge_mask_reg_512p3[11] <= 1'b1;
 		default: edge_mask_reg_512p3[11] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000101,
13'b11011000110,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100011000101,
13'b100011000110,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101011000101,
13'b101011000110,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110101,
13'b110010110110,
13'b111001000101,
13'b111001000110,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b1000001000101,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000001,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1010001000100,
13'b1010001000101,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010010001,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110001,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000001,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010010001,
13'b1011010010010,
13'b1011010010011,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001100001,
13'b1100001100010,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1100001110000,
13'b1100001110001,
13'b1100001110010,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100010000000,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010010001,
13'b1100010010010,
13'b1100010010011,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001010010,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001100001,
13'b1101001100010,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001110000,
13'b1101001110001,
13'b1101001110010,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101010000000,
13'b1101010000001,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010010001,
13'b1101010010010,
13'b1101010010011,
13'b1110001000011,
13'b1110001000100,
13'b1110001010010,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001100000,
13'b1110001100001,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001110000,
13'b1110001110001,
13'b1110001110010,
13'b1110001110011,
13'b1110001110100,
13'b1110001110101,
13'b1110010000000,
13'b1110010000001,
13'b1110010000010,
13'b1110010000011,
13'b1110010000100,
13'b1111001010011,
13'b1111001010100,
13'b1111001010101,
13'b1111001100000,
13'b1111001100001,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001100101,
13'b1111001110000,
13'b1111001110001,
13'b1111001110010,
13'b1111001110011,
13'b1111001110100,
13'b1111001110101,
13'b1111010000000,
13'b1111010000001,
13'b1111010000010: edge_mask_reg_512p3[12] <= 1'b1;
 		default: edge_mask_reg_512p3[12] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101111000,
13'b100101111001,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110001,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000000,
13'b100111000001,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101111000,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110001000,
13'b110110001001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110111000,
13'b111110111001,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111001000,
13'b111111001001,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111011000,
13'b111111011001,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111101000,
13'b1000110010011,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1001111000011,
13'b1001111010010,
13'b1001111010011,
13'b1001111100010,
13'b1001111100011: edge_mask_reg_512p3[13] <= 1'b1;
 		default: edge_mask_reg_512p3[13] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11110110111,
13'b11110111000,
13'b100110110111,
13'b100110111000,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100: edge_mask_reg_512p3[14] <= 1'b1;
 		default: edge_mask_reg_512p3[14] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101101000,
13'b10101101001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101111000,
13'b101101111001,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110001000,
13'b110110001001,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110011000,
13'b110110011001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001001,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111101000,
13'b111111101001,
13'b1000110010011,
13'b1000110010100,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001110100011,
13'b1001110100100,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1010111000100,
13'b1010111010100: edge_mask_reg_512p3[15] <= 1'b1;
 		default: edge_mask_reg_512p3[15] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101010111,
13'b101101011000,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111001000,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111011000,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111101000,
13'b111111101001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1010110000010,
13'b1010110000011,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111100000,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111110010,
13'b1010111110011,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011111000000,
13'b1011111000001,
13'b1100110100000,
13'b1100110100001: edge_mask_reg_512p3[16] <= 1'b1;
 		default: edge_mask_reg_512p3[16] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100110000111,
13'b100110001000,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101110000111,
13'b101110001000,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110010111,
13'b110110011000,
13'b110110100010,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111111000010,
13'b111111000011,
13'b111111000111,
13'b111111001000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010111,
13'b111111011000,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000111100010,
13'b1000111100011: edge_mask_reg_512p3[17] <= 1'b1;
 		default: edge_mask_reg_512p3[17] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000110,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110110,
13'b110000110111,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1001000010001,
13'b1001000010010,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011: edge_mask_reg_512p3[18] <= 1'b1;
 		default: edge_mask_reg_512p3[18] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000111,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100111,
13'b11011101000,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100111,
13'b100011101000,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100111,
13'b101011101000,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000001,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010111,
13'b110011011000,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001011000,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001101000,
13'b111001101001,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111011000000,
13'b111011000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010010000,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010100000,
13'b1000010100001,
13'b1000010100010,
13'b1000010110000,
13'b1000010110001,
13'b1000011000000,
13'b1001001000010,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001010000000,
13'b1001010000001,
13'b1001010000010,
13'b1001010010000,
13'b1001010010001,
13'b1001010010010,
13'b1001010100000,
13'b1001010100001,
13'b1001010110000,
13'b1001010110001,
13'b1010001100000,
13'b1010001100001,
13'b1010001110000,
13'b1010001110001,
13'b1010001110010,
13'b1010010000000,
13'b1010010000001,
13'b1010010010000,
13'b1010010010001,
13'b1010010100000,
13'b1010010100001,
13'b1011001110001: edge_mask_reg_512p3[19] <= 1'b1;
 		default: edge_mask_reg_512p3[19] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100111001,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b10001011010,
13'b10001011011,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110011,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110011,
13'b111011110100,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011011010,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110011,
13'b1000011110100,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1010010010111,
13'b1010010011000,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1011010011000,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011010111001,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011001001,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011011001,
13'b1011011100101,
13'b1011011100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100010111001,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011001001,
13'b1100011010111,
13'b1100011011000,
13'b1100011011001: edge_mask_reg_512p3[20] <= 1'b1;
 		default: edge_mask_reg_512p3[20] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100101001,
13'b100101010,
13'b100101011,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001011010,
13'b10001011011,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001011010,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011011010,
13'b1000011100011,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011100011,
13'b1001011100101,
13'b1001011100110,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011010111001,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011001001,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011011001,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100010111001,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011001001,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011011001: edge_mask_reg_512p3[21] <= 1'b1;
 		default: edge_mask_reg_512p3[21] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[22] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001001,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010001000,
13'b110010001001,
13'b110010011000,
13'b110010011001,
13'b111000010111,
13'b111000011000,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b1000000010111,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001011001,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001101001,
13'b1000001110111,
13'b1000001111000,
13'b1000001111001,
13'b1000010000111,
13'b1000010001000,
13'b1001000010111,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001000111000,
13'b1001001000110,
13'b1001001000111,
13'b1001001001000,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001101001,
13'b1001001110111,
13'b1001001111000,
13'b1001001111001,
13'b1001010000111,
13'b1001010001000,
13'b1010000010110,
13'b1010000010111,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010000111000,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001001000,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1010001100110,
13'b1010001100111,
13'b1010001101000,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1011001000101,
13'b1011001000110,
13'b1011001000111,
13'b1011001001000,
13'b1011001010101,
13'b1011001010110,
13'b1011001010111,
13'b1011001011000,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001100111,
13'b1011001101000,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011001110111,
13'b1011001111000,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010000111,
13'b1011010001000,
13'b1100000010101,
13'b1100000010110,
13'b1100000100101,
13'b1100000100110,
13'b1100000100111,
13'b1100000110100,
13'b1100000110101,
13'b1100000110110,
13'b1100000110111,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001000110,
13'b1100001000111,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001010111,
13'b1100001011000,
13'b1100001100100,
13'b1100001100101,
13'b1100001100110,
13'b1100001100111,
13'b1100001101000,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100001110111,
13'b1100001111000,
13'b1100010000100,
13'b1100010000101,
13'b1100010000110,
13'b1100010000111,
13'b1100010001000,
13'b1101000010101,
13'b1101000010110,
13'b1101000100101,
13'b1101000100110,
13'b1101000100111,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101000110110,
13'b1101000110111,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001000110,
13'b1101001000111,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001010110,
13'b1101001010111,
13'b1101001100100,
13'b1101001100101,
13'b1101001100110,
13'b1101001100111,
13'b1101001101000,
13'b1101001110100,
13'b1101001110101,
13'b1101001110110,
13'b1101001110111,
13'b1101001111000,
13'b1101010000100,
13'b1101010000101,
13'b1101010000110,
13'b1101010000111,
13'b1110000010101,
13'b1110000100101,
13'b1110000100110,
13'b1110000110011,
13'b1110000110100,
13'b1110000110101,
13'b1110000110110,
13'b1110000110111,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1110001000110,
13'b1110001000111,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001010110,
13'b1110001010111,
13'b1110001100100,
13'b1110001100101,
13'b1110001100110,
13'b1110001100111,
13'b1110001110100,
13'b1110001110101,
13'b1110001110110,
13'b1110001110111,
13'b1110010000100,
13'b1110010000101,
13'b1110010000111,
13'b1111000110011,
13'b1111000110100,
13'b1111000110101,
13'b1111000110110,
13'b1111001000011,
13'b1111001000100,
13'b1111001000101,
13'b1111001000110,
13'b1111001010100,
13'b1111001010101,
13'b1111001100100: edge_mask_reg_512p3[23] <= 1'b1;
 		default: edge_mask_reg_512p3[23] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100000,
13'b10010100001,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110000,
13'b10010110001,
13'b10010110010,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000000,
13'b10011000001,
13'b10011000010,
13'b10011000011,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010000,
13'b10011010010,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110010,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000000,
13'b11010000001,
13'b11010000010,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010000,
13'b11010010001,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100000,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110000,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000000,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010000,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100000,
13'b11011100001,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110000,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000000,
13'b11100000001,
13'b11100000010,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100101,
13'b11100100110,
13'b100000110101,
13'b100000110110,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100000,
13'b100001100001,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110000,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000000,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010000,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100000,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110000,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000000,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110000,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000000,
13'b100100000001,
13'b100100000010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100101,
13'b100100100110,
13'b101000110110,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000000,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110000,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000000,
13'b101100000001,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100101,
13'b101100100110,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010000,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110100000101,
13'b110100000110,
13'b110100010101,
13'b110100010110,
13'b111001010000,
13'b111001100000,
13'b111001100001,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110110,
13'b111001110111,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000000,
13'b111011000001,
13'b111011000010,
13'b111011000101,
13'b111011000110,
13'b111011010000,
13'b111011010001,
13'b111011010010,
13'b111011010101,
13'b111011010110,
13'b111011100000,
13'b111011100101,
13'b111011100110,
13'b1000001100000,
13'b1000001110000,
13'b1000001110001,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010010000,
13'b1000010010001,
13'b1000010010010,
13'b1000010100000,
13'b1000010100001,
13'b1000010110000,
13'b1000010110001,
13'b1001001110000,
13'b1001010000000: edge_mask_reg_512p3[24] <= 1'b1;
 		default: edge_mask_reg_512p3[24] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010111,
13'b11001011000,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010111,
13'b101001011000,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110001,
13'b110000110010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000100000,
13'b111000100001: edge_mask_reg_512p3[25] <= 1'b1;
 		default: edge_mask_reg_512p3[25] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100110101010,
13'b100110101011,
13'b100110110110,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110111000101,
13'b110111010100,
13'b110111010101,
13'b110111010110: edge_mask_reg_512p3[26] <= 1'b1;
 		default: edge_mask_reg_512p3[26] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100101,
13'b101100110,
13'b101100111,
13'b1101110101,
13'b1101110110,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101110000101,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111100000,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111110000,
13'b1010111110001,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111010000,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111100000,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111110000,
13'b1011111110001,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1100110110001,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111010000,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111100000,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111110000,
13'b1100111110001,
13'b1100111110010,
13'b1100111110011,
13'b1100111110100,
13'b1101111010000,
13'b1101111010001,
13'b1101111010010,
13'b1101111100000,
13'b1101111100001,
13'b1101111100010,
13'b1101111100011,
13'b1101111110000,
13'b1101111110001,
13'b1101111110010,
13'b1101111110011,
13'b1110111100000,
13'b1110111110000,
13'b1110111110001,
13'b1110111110010,
13'b1110111110011,
13'b1111111110000: edge_mask_reg_512p3[27] <= 1'b1;
 		default: edge_mask_reg_512p3[27] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[28] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[29] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100101,
13'b101100110,
13'b101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101110000101,
13'b101110000110,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111110110101,
13'b111110110110,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001110110100,
13'b1001110110101,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1010110110100,
13'b1010110110101,
13'b1010111000100,
13'b1010111000101,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1011110110100,
13'b1011110110101,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1101110110011,
13'b1101110110100,
13'b1101110110101,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111010011,
13'b1101111010100,
13'b1101111010101,
13'b1101111100011,
13'b1101111100100,
13'b1101111100101,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1110110110011,
13'b1110110110100,
13'b1110110110101,
13'b1110111000010,
13'b1110111000011,
13'b1110111000100,
13'b1110111000101,
13'b1110111010010,
13'b1110111010011,
13'b1110111010100,
13'b1110111010101,
13'b1110111100010,
13'b1110111100011,
13'b1110111100100,
13'b1110111100101,
13'b1110111110010,
13'b1110111110011,
13'b1110111110100,
13'b1110111110101,
13'b1111110110100,
13'b1111111000010,
13'b1111111000011,
13'b1111111000100,
13'b1111111000101,
13'b1111111010010,
13'b1111111010011,
13'b1111111010100,
13'b1111111010101,
13'b1111111100010,
13'b1111111100011,
13'b1111111100100,
13'b1111111100101,
13'b1111111110010,
13'b1111111110011,
13'b1111111110100,
13'b1111111110101: edge_mask_reg_512p3[30] <= 1'b1;
 		default: edge_mask_reg_512p3[30] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[31] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11110011010,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101110111010,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1000111101001,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1010111111000,
13'b1011111010110,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1011111110111,
13'b1011111111000,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110,
13'b1100111110111,
13'b1101111110100,
13'b1101111110101: edge_mask_reg_512p3[32] <= 1'b1;
 		default: edge_mask_reg_512p3[32] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b100011101000,
13'b100011101001,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b110011111000,
13'b110011111001,
13'b110100001000,
13'b110100001001,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110011000,
13'b110110011001,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000101,
13'b111110000110,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000100,
13'b1001110000101,
13'b1010100010100,
13'b1010100010101,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000010,
13'b1010110000100,
13'b1010110000101,
13'b1011100010100,
13'b1011100010101,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1100100100011,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100100110101,
13'b1100100110110,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1101100100011,
13'b1101100100100,
13'b1101100100101,
13'b1101100110010,
13'b1101100110011,
13'b1101100110100,
13'b1101100110101,
13'b1101100110110,
13'b1101101000010,
13'b1101101000011,
13'b1101101000100,
13'b1101101000101,
13'b1101101000110,
13'b1101101010010,
13'b1101101010011,
13'b1101101010100,
13'b1101101010101,
13'b1101101100010,
13'b1101101100011,
13'b1110100100011,
13'b1110100100100,
13'b1110100110010,
13'b1110100110011,
13'b1110100110100,
13'b1110101000010,
13'b1110101000011,
13'b1110101000100,
13'b1110101010011,
13'b1111100110011,
13'b1111101000011,
13'b1111101000100: edge_mask_reg_512p3[33] <= 1'b1;
 		default: edge_mask_reg_512p3[33] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[34] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[35] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b100111001010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101011010,
13'b1000101101000,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101111000,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1000110001000,
13'b1000110001001,
13'b1000110001010,
13'b1000110001011,
13'b1000110011000,
13'b1000110011001,
13'b1001101011000,
13'b1001101011001,
13'b1001101011010,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101101010,
13'b1001101111000,
13'b1001101111001,
13'b1001101111010,
13'b1001101111011,
13'b1001110001000,
13'b1001110001001,
13'b1001110001010,
13'b1001110001011,
13'b1001110011000,
13'b1001110011001,
13'b1010101011000,
13'b1010101011001,
13'b1010101011010,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101101010,
13'b1010101111000,
13'b1010101111001,
13'b1010101111010,
13'b1010101111011,
13'b1010110001000,
13'b1010110001001,
13'b1010110001010,
13'b1010110001011,
13'b1010110011000,
13'b1010110011001,
13'b1011101010111,
13'b1011101011000,
13'b1011101011001,
13'b1011101011010,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1011101101010,
13'b1011101110111,
13'b1011101111000,
13'b1011101111001,
13'b1011101111010,
13'b1011101111011,
13'b1011110000111,
13'b1011110001000,
13'b1011110001001,
13'b1011110001010,
13'b1011110011000,
13'b1011110011001,
13'b1100101010111,
13'b1100101011000,
13'b1100101011001,
13'b1100101011010,
13'b1100101100111,
13'b1100101101000,
13'b1100101101001,
13'b1100101101010,
13'b1100101101011,
13'b1100101110111,
13'b1100101111000,
13'b1100101111001,
13'b1100101111010,
13'b1100101111011,
13'b1100110000111,
13'b1100110001000,
13'b1100110001001,
13'b1100110001010,
13'b1100110001011,
13'b1100110011000,
13'b1101101010111,
13'b1101101011000,
13'b1101101011001,
13'b1101101011010,
13'b1101101100111,
13'b1101101101000,
13'b1101101101001,
13'b1101101101010,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101101111001,
13'b1101101111010,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1101110001001,
13'b1101110001010,
13'b1101110011000,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101101001,
13'b1110101101010,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110101111001,
13'b1110101111010,
13'b1110110000101,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110001001,
13'b1110110001010,
13'b1111101100110,
13'b1111101100111,
13'b1111101101000,
13'b1111101101001,
13'b1111101110101,
13'b1111101110110,
13'b1111101110111,
13'b1111101111000,
13'b1111101111001,
13'b1111110000101,
13'b1111110000110,
13'b1111110000111,
13'b1111110001000: edge_mask_reg_512p3[36] <= 1'b1;
 		default: edge_mask_reg_512p3[36] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11010101,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110101,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100000,
13'b100100001,
13'b100100110,
13'b100100111,
13'b100110000,
13'b100110001,
13'b100110110,
13'b100110111,
13'b101000000,
13'b101000001,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000000,
13'b1100000001,
13'b1100000010,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010000,
13'b1100010001,
13'b1100010010,
13'b1100010011,
13'b1100010100,
13'b1100010110,
13'b1100010111,
13'b1100100000,
13'b1100100001,
13'b1100100010,
13'b1100100011,
13'b1100100100,
13'b1100110000,
13'b1100110001,
13'b1100110010,
13'b1100110011,
13'b1101000000,
13'b1101000001,
13'b1101000010,
13'b1101000011,
13'b1101010000,
13'b1101010001,
13'b1101010110,
13'b1101010111,
13'b1101100000,
13'b1101100001,
13'b1101100010,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110000,
13'b10011110001,
13'b10011110010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000000,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010000,
13'b10100010001,
13'b10100010010,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100000,
13'b10100100001,
13'b10100100010,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110000,
13'b10100110001,
13'b10100110010,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000000,
13'b10101000001,
13'b10101000010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010000,
13'b10101010001,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100000,
13'b10101100001,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110000,
13'b10101110001,
13'b10101110010,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b11011100110,
13'b11011100111,
13'b11011110000,
13'b11011110001,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000000,
13'b11100000001,
13'b11100000010,
13'b11100000011,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010000,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100000,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110000,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000000,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010000,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010000,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100000,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b110011110110,
13'b110011110111,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111101000101,
13'b111101000110,
13'b111101000111: edge_mask_reg_512p3[37] <= 1'b1;
 		default: edge_mask_reg_512p3[37] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101100111,
13'b101101000,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b110100011000,
13'b110100011001,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b1000100100011,
13'b1000100100100,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000011,
13'b1001110000100,
13'b1010100110001,
13'b1010100110010,
13'b1010101000001,
13'b1010101000010,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101110010,
13'b1010101110011,
13'b1011101000001,
13'b1011101000010,
13'b1011101010001,
13'b1011101010010,
13'b1011101100010: edge_mask_reg_512p3[38] <= 1'b1;
 		default: edge_mask_reg_512p3[38] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110100011000,
13'b110100011001,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101011000,
13'b111101011001,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101101000,
13'b111101101001,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101111000,
13'b111101111001,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110001000,
13'b111110001001,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110011000,
13'b111110011001,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110101000,
13'b111110101001,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110111000,
13'b111110111001,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111001000,
13'b111111001001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110100000,
13'b1001110100001,
13'b1010100110001,
13'b1010100110010,
13'b1010101000001,
13'b1010101000010,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101100001,
13'b1010101100010,
13'b1010101110001,
13'b1010101110010,
13'b1010110000001,
13'b1011101000001,
13'b1011101000010,
13'b1011101010001,
13'b1011101010010,
13'b1011101100001: edge_mask_reg_512p3[39] <= 1'b1;
 		default: edge_mask_reg_512p3[39] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100110,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b101011011001,
13'b101011011010,
13'b101011100101,
13'b101011100110,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101111000,
13'b110101111001,
13'b110110001000,
13'b110110001001,
13'b111011100100,
13'b111011100101,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110011,
13'b1000101110100,
13'b1001011110010,
13'b1001011110011,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010010,
13'b1010100010011,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1011100000011,
13'b1011100010010,
13'b1011100010011,
13'b1011100110010,
13'b1011101000001,
13'b1011101000010,
13'b1011101010001,
13'b1011101010010: edge_mask_reg_512p3[40] <= 1'b1;
 		default: edge_mask_reg_512p3[40] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101001000,
13'b11101001001,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100101001001,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101101000,
13'b110101101001,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111001000,
13'b110111001001,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1100110000010,
13'b1100110000011,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1101110010010,
13'b1101110010011,
13'b1101110100010,
13'b1101110100011: edge_mask_reg_512p3[41] <= 1'b1;
 		default: edge_mask_reg_512p3[41] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101001000,
13'b11101001001,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100101001001,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b101111011011,
13'b110101101000,
13'b110101101001,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111100100,
13'b1001111100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111010010,
13'b1010111010011,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110110010,
13'b1011110110011,
13'b1011111000010,
13'b1011111000011,
13'b1100110000010,
13'b1100110010010,
13'b1100110010011,
13'b1100110100010,
13'b1100110100011,
13'b1100110110010,
13'b1101110010010,
13'b1101110100010: edge_mask_reg_512p3[42] <= 1'b1;
 		default: edge_mask_reg_512p3[42] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101001000,
13'b11101001001,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101001001,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1100110000001,
13'b1100110000010,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110100000,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110110000,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1101110010010,
13'b1101110100001,
13'b1101110100010,
13'b1101110110001: edge_mask_reg_512p3[43] <= 1'b1;
 		default: edge_mask_reg_512p3[43] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10011101000,
13'b10011101001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101011111001,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110100001001,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111001000,
13'b110111001001,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1011101000010,
13'b1011101010010,
13'b1011101010011,
13'b1011101100010,
13'b1011101100011,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1100101100010,
13'b1100101110010,
13'b1100110000010,
13'b1100110000011,
13'b1100110010010,
13'b1100110010011,
13'b1100110100010,
13'b1100110100011,
13'b1101110010010: edge_mask_reg_512p3[44] <= 1'b1;
 		default: edge_mask_reg_512p3[44] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b1001100110,
13'b1001100111,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000111,
13'b11011001000,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110000,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000000,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000111,
13'b100011001000,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000111,
13'b101011001000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100001,
13'b110010100010,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110111,
13'b110010111000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110110,
13'b111000110111,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100111,
13'b111001101000,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110111,
13'b111001111000,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000111,
13'b111010001000,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b1000000100001,
13'b1000000100010,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100: edge_mask_reg_512p3[45] <= 1'b1;
 		default: edge_mask_reg_512p3[45] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100010,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110001,
13'b101001110010,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000001,
13'b101010000010,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010001,
13'b101010010010,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110010,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100001,
13'b110010100100,
13'b110010100101,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001001,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010100001,
13'b111010100010,
13'b111010100100,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000010111,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010010011,
13'b1010010010100,
13'b1011000000100,
13'b1011000000101,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000010110,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001110011,
13'b1011001110100,
13'b1100000010100,
13'b1100000010101,
13'b1100000100100,
13'b1100000100101,
13'b1100000110100,
13'b1100000110101,
13'b1100001000100,
13'b1100001000101: edge_mask_reg_512p3[46] <= 1'b1;
 		default: edge_mask_reg_512p3[46] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1010100101,
13'b1010100110,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b11010110101,
13'b11010110110,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b100010110101,
13'b100010110110,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b111011100000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110110,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000110,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010110,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100110,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110110,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1010011100000,
13'b1010011100001,
13'b1010011110000,
13'b1010011110001,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1011100000000,
13'b1011100000001,
13'b1011100010000,
13'b1011100010001,
13'b1011100100000,
13'b1011100100001,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101100000,
13'b1011101100001,
13'b1011101100010,
13'b1100100000000,
13'b1100100010000,
13'b1100100100000,
13'b1100100110000,
13'b1100100110001,
13'b1100101000000,
13'b1100101000001,
13'b1100101010000,
13'b1100101010001,
13'b1100101100000,
13'b1100101100001,
13'b1101100100000,
13'b1101100110000,
13'b1101101000000,
13'b1101101000001,
13'b1101101010000,
13'b1101101010001,
13'b1101101100000,
13'b1110100110000,
13'b1110101000000,
13'b1110101010000: edge_mask_reg_512p3[47] <= 1'b1;
 		default: edge_mask_reg_512p3[47] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100101000,
13'b100101001,
13'b100101010,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b11001001010,
13'b11001001011,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b101001110111,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110101,
13'b101011111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110100,
13'b110011110101,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011100100,
13'b111011100101,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000011,
13'b1010011000100,
13'b1011010010100,
13'b1011010100100,
13'b1011010110100: edge_mask_reg_512p3[48] <= 1'b1;
 		default: edge_mask_reg_512p3[48] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b100111010,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b11001001010,
13'b11001001011,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b101001110111,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1011010010100,
13'b1011010010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1100010100100,
13'b1100010110100,
13'b1100010110101,
13'b1100011000100,
13'b1100011000101,
13'b1100011010100,
13'b1100011010101,
13'b1101011000100,
13'b1101011010100: edge_mask_reg_512p3[49] <= 1'b1;
 		default: edge_mask_reg_512p3[49] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101010,
13'b11001001010,
13'b11001001011,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101001110111,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100100,
13'b1001100100101,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1011010010100,
13'b1011010100100,
13'b1011010110011,
13'b1011010110100,
13'b1011011000011,
13'b1011011000100,
13'b1011011010011,
13'b1011011010100,
13'b1011011100011,
13'b1011011100100,
13'b1011011110011,
13'b1011011110100,
13'b1011100000011,
13'b1011100000100: edge_mask_reg_512p3[50] <= 1'b1;
 		default: edge_mask_reg_512p3[50] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101011001,
13'b1101011010,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11001001010,
13'b11001001011,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101011010,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b101001110111,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010101,
13'b1011010010100,
13'b1011010100100,
13'b1011010100101,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011100011,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011110011,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1100010110100,
13'b1100011000100,
13'b1100011010011,
13'b1100011010100,
13'b1100011100011,
13'b1100011100100,
13'b1100011110011,
13'b1100011110100,
13'b1100011110101,
13'b1100100000011,
13'b1100100000100,
13'b1100100000101,
13'b1101011100100,
13'b1101011110100,
13'b1101100000100: edge_mask_reg_512p3[51] <= 1'b1;
 		default: edge_mask_reg_512p3[51] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100111000,
13'b101100111001,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110100,
13'b1000110110101,
13'b1001101010001,
13'b1001101010011,
13'b1001101010100,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110110100,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110100011,
13'b1010110100100,
13'b1010110110011,
13'b1010110110100,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110100011,
13'b1011110100100,
13'b1100110000001,
13'b1100110000010: edge_mask_reg_512p3[52] <= 1'b1;
 		default: edge_mask_reg_512p3[52] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[53] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[54] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11011101,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11101101,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b11111101,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100001101,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101101011,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011011101,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011101101,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1011111101,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100001101,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101011,
13'b10001101010,
13'b10001101011,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011011101,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011101101,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10011111101,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b100010001010,
13'b100010001011,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011010,
13'b100100011011,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b110010100111,
13'b110010101000,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011011011,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011011010,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1000011101010,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000011111010,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100001010,
13'b1001010100110,
13'b1001010100111,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011001010,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011011010,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011101001,
13'b1001011101010,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001011111001,
13'b1001011111010,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100001010,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1010011011010,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011101001,
13'b1010011101010,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010011111001,
13'b1010011111010,
13'b1010100000111,
13'b1010100001000,
13'b1010100001001,
13'b1010100001010,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011001001,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011011001,
13'b1011011011010,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011101000,
13'b1011011101001,
13'b1011011101010,
13'b1011011110110,
13'b1011011110111,
13'b1011011111000,
13'b1011011111001,
13'b1011011111010,
13'b1011100001000,
13'b1011100001001,
13'b1100011000101,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1100011101001,
13'b1100011110110,
13'b1100011110111,
13'b1100011111000,
13'b1100011111001,
13'b1101011010110,
13'b1101011010111,
13'b1101011100110,
13'b1101011100111,
13'b1101011101000,
13'b1101011110110,
13'b1101011110111,
13'b1101011111000: edge_mask_reg_512p3[55] <= 1'b1;
 		default: edge_mask_reg_512p3[55] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10011110110,
13'b10011110111,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101100000110,
13'b101100000111,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110111,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110110,
13'b111110110111,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111010000,
13'b1000100100001,
13'b1000100100010,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1001100110001,
13'b1001100110010,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110100001,
13'b1001110100010,
13'b1001110110001,
13'b1001110110010,
13'b1010101000001,
13'b1010101000010,
13'b1010101010001,
13'b1010101010010,
13'b1010101100001,
13'b1010101100010,
13'b1010101110001,
13'b1010101110010,
13'b1010110000001,
13'b1010110000010,
13'b1010110010001: edge_mask_reg_512p3[56] <= 1'b1;
 		default: edge_mask_reg_512p3[56] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111100,
13'b101001011,
13'b101001100,
13'b101011011,
13'b101011100,
13'b101011101,
13'b101101010,
13'b101101011,
13'b101101100,
13'b101101101,
13'b1101111011,
13'b1101111100,
13'b1110001011,
13'b1110001100,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b1110011101,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b10110101010,
13'b11110011001,
13'b11110101000,
13'b11110101001,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110100101,
13'b110110100110,
13'b110110101000,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110110101,
13'b111110110110,
13'b111111000101,
13'b111111000110,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000111100101: edge_mask_reg_512p3[57] <= 1'b1;
 		default: edge_mask_reg_512p3[57] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101001,
13'b10101101010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101001,
13'b11101101010,
13'b100001011000,
13'b100001011001,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010001,
13'b100010010010,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110101,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110001110011,
13'b110001110100,
13'b110001111000,
13'b110001111001,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010001000,
13'b110010001001,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011001,
13'b110010011010,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b1000010000011,
13'b1000010000100,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1001010100011,
13'b1001010100100,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110100,
13'b1001100110101,
13'b1010011000100,
13'b1010011010001,
13'b1010011010010,
13'b1010011010100,
13'b1010011010101,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110100,
13'b1010100110101,
13'b1011011110010,
13'b1011011110011,
13'b1011011110101,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1100100010010: edge_mask_reg_512p3[58] <= 1'b1;
 		default: edge_mask_reg_512p3[58] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100001,
13'b100001100010,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110001,
13'b100001110010,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000001,
13'b100010000010,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b101000100101,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110001,
13'b101000110010,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b110000100101,
13'b110000101000,
13'b110000101001,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001000,
13'b110011001001,
13'b110011010011,
13'b110011010100,
13'b110011011001,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111011000011,
13'b111011000100,
13'b111011010011,
13'b111011010100,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010110011,
13'b1000010110100,
13'b1001000110011,
13'b1001000110100,
13'b1001001000011,
13'b1001001000100,
13'b1001001010011,
13'b1001001010100,
13'b1001001100011,
13'b1001001100100: edge_mask_reg_512p3[59] <= 1'b1;
 		default: edge_mask_reg_512p3[59] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b100001011000,
13'b100001011001,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010001,
13'b100010010010,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110101,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b110001110011,
13'b110001110100,
13'b110001111000,
13'b110001111001,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010001001,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011001,
13'b110010011010,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101010,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000111,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000101,
13'b1000010000011,
13'b1000010000100,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000101,
13'b1001010010100,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000101,
13'b1010010110100,
13'b1010010110101,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100101: edge_mask_reg_512p3[60] <= 1'b1;
 		default: edge_mask_reg_512p3[60] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[61] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110111,
13'b1011111000,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b101000101001,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b110000111001,
13'b110001001000,
13'b110001001001,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110111,
13'b111010111000,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001101001,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000001111001,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010001001,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110111,
13'b1000010111000,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001001111001,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010001001,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110111,
13'b1001010111000,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1010001100110,
13'b1010001100111,
13'b1010001101000,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110111,
13'b1010010111000,
13'b1011001010101,
13'b1011001010110,
13'b1011001010111,
13'b1011001100101,
13'b1011001100110,
13'b1011001100111,
13'b1011001101000,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011001110111,
13'b1011001111000,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010000111,
13'b1011010001000,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1100001010101,
13'b1100001010110,
13'b1100001010111,
13'b1100001100101,
13'b1100001100110,
13'b1100001100111,
13'b1100001101000,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100001110111,
13'b1100001111000,
13'b1100010000100,
13'b1100010000101,
13'b1100010000110,
13'b1100010000111,
13'b1100010001000,
13'b1100010010100,
13'b1100010010101,
13'b1100010010110,
13'b1100010010111,
13'b1100010011000,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1101001010110,
13'b1101001010111,
13'b1101001100100,
13'b1101001100101,
13'b1101001100110,
13'b1101001100111,
13'b1101001101000,
13'b1101001110100,
13'b1101001110101,
13'b1101001110110,
13'b1101001110111,
13'b1101001111000,
13'b1101010000100,
13'b1101010000101,
13'b1101010000110,
13'b1101010000111,
13'b1101010001000,
13'b1101010010100,
13'b1101010010101,
13'b1101010010110,
13'b1101010010111,
13'b1101010011000,
13'b1101010100100,
13'b1101010100101,
13'b1101010100110,
13'b1101010100111,
13'b1101010101000,
13'b1101010110100,
13'b1101010110101,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000100,
13'b1101011000101,
13'b1110001100110,
13'b1110001100111,
13'b1110001110100,
13'b1110001110101,
13'b1110001110110,
13'b1110001110111,
13'b1110010000100,
13'b1110010000101,
13'b1110010000110,
13'b1110010000111,
13'b1110010001000,
13'b1110010010100,
13'b1110010010101,
13'b1110010010110,
13'b1110010010111,
13'b1110010011000,
13'b1110010100100,
13'b1110010100101,
13'b1110010100110,
13'b1110010100111,
13'b1110010101000,
13'b1110010110100,
13'b1110010110101,
13'b1110010110110,
13'b1110010110111,
13'b1110011000100,
13'b1110011000101,
13'b1111010010100,
13'b1111010010101,
13'b1111010010110,
13'b1111010010111,
13'b1111010100100,
13'b1111010100101,
13'b1111010100110,
13'b1111010100111,
13'b1111010110100,
13'b1111010110101,
13'b1111010110111: edge_mask_reg_512p3[62] <= 1'b1;
 		default: edge_mask_reg_512p3[62] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000110,
13'b11000111,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110110,
13'b100110111,
13'b101000110,
13'b101000111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110110,
13'b1100110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110110,
13'b10100110111,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110110,
13'b11100110111,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110110,
13'b100100110111,
13'b101010000110,
13'b101010000111,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110110,
13'b101100110111,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100110,
13'b110100100111,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1011010110010,
13'b1011010110011,
13'b1011010110100,
13'b1011011000001,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011010100,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000010,
13'b1011100000011,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100011000001,
13'b1100011000010,
13'b1100011000011,
13'b1100011000100,
13'b1100011010000,
13'b1100011010001,
13'b1100011010010,
13'b1100011010011,
13'b1100011010100,
13'b1100011100000,
13'b1100011100001,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011110000,
13'b1100011110001,
13'b1100011110010,
13'b1100011110011,
13'b1100100000010,
13'b1100100000011,
13'b1101010110010,
13'b1101010110011,
13'b1101011000001,
13'b1101011000010,
13'b1101011000011,
13'b1101011000100,
13'b1101011010000,
13'b1101011010001,
13'b1101011010010,
13'b1101011010011,
13'b1101011010100,
13'b1101011100000,
13'b1101011100001,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011110000,
13'b1101011110001,
13'b1101011110010,
13'b1101011110011,
13'b1110011000000,
13'b1110011000001,
13'b1110011000010,
13'b1110011000011,
13'b1110011010000,
13'b1110011010001,
13'b1110011010010,
13'b1110011010011,
13'b1110011100000,
13'b1110011100001,
13'b1110011100010,
13'b1110011110000,
13'b1110011110001,
13'b1111011000000,
13'b1111011000001,
13'b1111011000010,
13'b1111011010000,
13'b1111011010001,
13'b1111011010010,
13'b1111011100001,
13'b1111011100010,
13'b1111011110001: edge_mask_reg_512p3[63] <= 1'b1;
 		default: edge_mask_reg_512p3[63] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011001001,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001001011,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101001,
13'b101010101010,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b111000010110,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010010,
13'b111001010011,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b1000000010101,
13'b1000000010110,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1001000010101,
13'b1001000010110,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1011000010100,
13'b1011000010101,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110101,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000110010,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100000110110,
13'b1100001000010,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001010100,
13'b1100001010101: edge_mask_reg_512p3[64] <= 1'b1;
 		default: edge_mask_reg_512p3[64] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010100,
13'b100010101,
13'b100010110,
13'b100100100,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110100,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000100,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010100,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100100,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10100100100,
13'b10100100101,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000011,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010011,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100011,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101100110100,
13'b101100110101,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b110101000100,
13'b110101000101,
13'b110101010000,
13'b110101010001,
13'b110101010100,
13'b110101010101,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b111101100000,
13'b111101100001,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000101,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b1000101100000,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1001101110000,
13'b1001110000000,
13'b1001110000001,
13'b1001110010000,
13'b1001110010001,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001111000000,
13'b1001111000001,
13'b1010110000000,
13'b1010110000001,
13'b1010110010000,
13'b1010110010001,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010111000000,
13'b1011110010000,
13'b1011110100000,
13'b1011110100001,
13'b1011110110000,
13'b1011110110001: edge_mask_reg_512p3[65] <= 1'b1;
 		default: edge_mask_reg_512p3[65] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[66] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100111001,
13'b100111010,
13'b100111011,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010000010,
13'b1010000011,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010010010,
13'b1010010011,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010100010,
13'b1010100011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010110010,
13'b1010110011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111010,
13'b1100111011,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001110010,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010000010,
13'b10010000011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010010010,
13'b10010010011,
13'b10010010100,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010100010,
13'b10010100011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010110010,
13'b10010110011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011000010,
13'b10011000011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101010,
13'b10100101011,
13'b10100111010,
13'b10100111011,
13'b11001001001,
13'b11001001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110010,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000010,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011000010,
13'b11011000011,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101010,
13'b11100101011,
13'b100001001001,
13'b100001001010,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100100,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b101001100101,
13'b101001101001,
13'b101001101010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111001,
13'b101001111010,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b111001110100,
13'b111001110101,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b1000010000100,
13'b1000010000101,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1010010100110,
13'b1010010100111,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000110,
13'b1010011000111,
13'b1010011010110,
13'b1010011010111: edge_mask_reg_512p3[67] <= 1'b1;
 		default: edge_mask_reg_512p3[67] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b1001100100,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110100,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000100,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b11001000011,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110101,
13'b11010110110,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010110101,
13'b100010110110,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100101,
13'b110010100110,
13'b111000010000,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000010,
13'b111010000011,
13'b1000000010000,
13'b1000000010001,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000010000010,
13'b1000010000011,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001010000001,
13'b1001010000010,
13'b1001010000011,
13'b1010000100000,
13'b1010000100001,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001110000,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001010000,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001100000,
13'b1011001100001,
13'b1011001100010,
13'b1011001110000,
13'b1011001110001,
13'b1011001110010,
13'b1011001110011,
13'b1011010000001,
13'b1011010000010,
13'b1100001000001,
13'b1100001000010,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001100000,
13'b1100001100001,
13'b1100001100010,
13'b1100001110001,
13'b1100001110010,
13'b1100010000001,
13'b1100010000010: edge_mask_reg_512p3[68] <= 1'b1;
 		default: edge_mask_reg_512p3[68] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[69] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[70] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[71] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[72] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11010110,
13'b11010111,
13'b11100110,
13'b11100111,
13'b11110110,
13'b11110111,
13'b100000110,
13'b100000111,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011100110,
13'b1011100111,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10011100110,
13'b10011100111,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101011110110,
13'b101011110111,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010010,
13'b101100010011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010110,
13'b101111010111,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100110,
13'b111100100111,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110001,
13'b1000110110010,
13'b1001100100001,
13'b1001100100010,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110001,
13'b1001110110010,
13'b1010101000001,
13'b1010101000010,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1011101100000,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1100101110000,
13'b1100110000000,
13'b1100110000001,
13'b1100110010000: edge_mask_reg_512p3[73] <= 1'b1;
 		default: edge_mask_reg_512p3[73] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100010101,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101110111,
13'b1110010110,
13'b1110010111,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11100100101,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010110,
13'b101111010111,
13'b110101000001,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110001,
13'b1000110110010,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110001,
13'b1001110110010,
13'b1010101100001,
13'b1010101100010,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1100110000000,
13'b1100110000001,
13'b1100110010000: edge_mask_reg_512p3[74] <= 1'b1;
 		default: edge_mask_reg_512p3[74] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100110,
13'b100100111,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100110110,
13'b1100110111,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101101000110,
13'b101101000111,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100101,
13'b111111100110,
13'b1000101100011,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111100000,
13'b1000111100001,
13'b1001101100011,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111010000,
13'b1001111010001,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010111000001,
13'b1010111000010,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1100110000000,
13'b1100110000001,
13'b1100110010000: edge_mask_reg_512p3[75] <= 1'b1;
 		default: edge_mask_reg_512p3[75] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100110,
13'b100100111,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100110110,
13'b1100110111,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101000110,
13'b101101000111,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b1000101100011,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1001101100011,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111010010,
13'b1011111010011,
13'b1100110000000,
13'b1100110000001,
13'b1100110010000,
13'b1100110010001,
13'b1100110100000,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110110000,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1101110010000,
13'b1101110100000,
13'b1101110100001,
13'b1101110110000,
13'b1101110110001: edge_mask_reg_512p3[76] <= 1'b1;
 		default: edge_mask_reg_512p3[76] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100110,
13'b100100111,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100110110,
13'b1100110111,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101000110,
13'b101101000111,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b1000101100011,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001101100011,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1100110000000,
13'b1100110000001,
13'b1100110010000,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110100000,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1100110110000,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1101110000000,
13'b1101110010000,
13'b1101110010001,
13'b1101110010010,
13'b1101110100000,
13'b1101110100001,
13'b1101110100010,
13'b1101110100011,
13'b1101110110000,
13'b1101110110001,
13'b1101110110010,
13'b1101110110011,
13'b1101110110100,
13'b1101111000001,
13'b1101111000010,
13'b1101111000011,
13'b1101111000100,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1110110010001,
13'b1110110100001,
13'b1110110100010,
13'b1110110110001,
13'b1110110110010,
13'b1110110110011,
13'b1110111000001,
13'b1110111000010,
13'b1110111000011,
13'b1110111000100,
13'b1110111010010,
13'b1110111010011,
13'b1110111010100,
13'b1111110110001,
13'b1111110110010,
13'b1111110110011,
13'b1111111000010,
13'b1111111000011,
13'b1111111000100,
13'b1111111010010,
13'b1111111010011: edge_mask_reg_512p3[77] <= 1'b1;
 		default: edge_mask_reg_512p3[77] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b1001100010,
13'b1001100011,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001110010,
13'b1001110011,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011011000,
13'b1011011001,
13'b10001010010,
13'b10001010011,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100010,
13'b10001100011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001110010,
13'b10001110011,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000010,
13'b10010000011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010010,
13'b10010010011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b11001000010,
13'b11001000011,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001010010,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100010,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110010,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000010,
13'b11010000011,
13'b11010000100,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011001,
13'b11011011010,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010010,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110010,
13'b101010110011,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001001,
13'b101011001010,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000101000,
13'b110000101001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000101000,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000111000,
13'b111000111001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001001000,
13'b111001001001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b1000000110011,
13'b1000001000011,
13'b1000001000100,
13'b1000001010011,
13'b1000001010100,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1001001110011,
13'b1001001110100,
13'b1001010000011,
13'b1001010000100,
13'b1001010010011,
13'b1001010010100: edge_mask_reg_512p3[78] <= 1'b1;
 		default: edge_mask_reg_512p3[78] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11010110,
13'b11010111,
13'b11100110,
13'b11100111,
13'b11110110,
13'b11110111,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011100110,
13'b1011100111,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011100110,
13'b10011100111,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101011110110,
13'b101011110111,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010010,
13'b101100010011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010110,
13'b110111010111,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100110,
13'b111100100111,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1001100100001,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110110001,
13'b1010110110010,
13'b1011101110000,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010: edge_mask_reg_512p3[79] <= 1'b1;
 		default: edge_mask_reg_512p3[79] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100010101,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110110,
13'b1101110111,
13'b1110010110,
13'b1110010111,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11100100101,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110101000001,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010110,
13'b110111010111,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100101,
13'b111101100110,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b1000101010000,
13'b1000101010001,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010: edge_mask_reg_512p3[80] <= 1'b1;
 		default: edge_mask_reg_512p3[80] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10100000101,
13'b10100000110,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101100010101,
13'b101100010110,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010110,
13'b110111010111,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000101,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b1000100110000,
13'b1000100110001,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1001101000000,
13'b1001101000001,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110110001,
13'b1010110110010,
13'b1011101110000,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010: edge_mask_reg_512p3[81] <= 1'b1;
 		default: edge_mask_reg_512p3[81] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100101000110,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110101010110,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100101,
13'b111111100110,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111100000,
13'b1000111100001,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111010000,
13'b1001111010001,
13'b1010101110001,
13'b1010101110010,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010: edge_mask_reg_512p3[82] <= 1'b1;
 		default: edge_mask_reg_512p3[82] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101000110,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101010110,
13'b110101010111,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1010101110001,
13'b1010101110010,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111010010,
13'b1011111010011,
13'b1100110000000,
13'b1100110010000,
13'b1100110010001,
13'b1100110100000,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110110000,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1101110100000,
13'b1101110100001,
13'b1101110110000,
13'b1101110110001: edge_mask_reg_512p3[83] <= 1'b1;
 		default: edge_mask_reg_512p3[83] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101101000110,
13'b101101000111,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010110,
13'b110111010111,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b1000101100011,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1001101100011,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110110001,
13'b1010110110010,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1100110000000,
13'b1100110000001,
13'b1100110010000: edge_mask_reg_512p3[84] <= 1'b1;
 		default: edge_mask_reg_512p3[84] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[85] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110011011001,
13'b110011011010,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b1000011011001,
13'b1000011011010,
13'b1000011011011,
13'b1000011101001,
13'b1000011101010,
13'b1000011101011,
13'b1000011111001,
13'b1000011111010,
13'b1000011111011,
13'b1000100001001,
13'b1000100001010,
13'b1000100001011,
13'b1000100011001,
13'b1000100011010,
13'b1000100011011,
13'b1000100101001,
13'b1000100101010,
13'b1000100101011,
13'b1000100111001,
13'b1000100111010,
13'b1000100111011,
13'b1000101001011,
13'b1001011011001,
13'b1001011011010,
13'b1001011011011,
13'b1001011101001,
13'b1001011101010,
13'b1001011101011,
13'b1001011111001,
13'b1001011111010,
13'b1001011111011,
13'b1001100001001,
13'b1001100001010,
13'b1001100001011,
13'b1001100011001,
13'b1001100011010,
13'b1001100011011,
13'b1001100101001,
13'b1001100101010,
13'b1001100101011,
13'b1001100111010,
13'b1001100111011,
13'b1001101001011,
13'b1010011011010,
13'b1010011011011,
13'b1010011101010,
13'b1010011101011,
13'b1010011111010,
13'b1010011111011,
13'b1010011111100,
13'b1010100001001,
13'b1010100001010,
13'b1010100001011,
13'b1010100001100,
13'b1010100011001,
13'b1010100011010,
13'b1010100011011,
13'b1010100011100,
13'b1010100101010,
13'b1010100101011,
13'b1010100101100,
13'b1010100111010,
13'b1010100111011,
13'b1010100111100,
13'b1010101001011,
13'b1011011011010,
13'b1011011011011,
13'b1011011101010,
13'b1011011101011,
13'b1011011101100,
13'b1011011111010,
13'b1011011111011,
13'b1011011111100,
13'b1011100001010,
13'b1011100001011,
13'b1011100001100,
13'b1011100011010,
13'b1011100011011,
13'b1011100011100,
13'b1011100101010,
13'b1011100101011,
13'b1011100101100,
13'b1011100111010,
13'b1011100111011,
13'b1011100111100,
13'b1011101001011,
13'b1011101001100,
13'b1100011011010,
13'b1100011011011,
13'b1100011011100,
13'b1100011101010,
13'b1100011101011,
13'b1100011101100,
13'b1100011111010,
13'b1100011111011,
13'b1100011111100,
13'b1100100001010,
13'b1100100001011,
13'b1100100001100,
13'b1100100011010,
13'b1100100011011,
13'b1100100011100,
13'b1100100101010,
13'b1100100101011,
13'b1100100101100,
13'b1100100111010,
13'b1100100111011,
13'b1100100111100,
13'b1100101001011,
13'b1100101001100,
13'b1101011011010,
13'b1101011011011,
13'b1101011011100,
13'b1101011101010,
13'b1101011101011,
13'b1101011101100,
13'b1101011111010,
13'b1101011111011,
13'b1101011111100,
13'b1101100001010,
13'b1101100001011,
13'b1101100001100,
13'b1101100011010,
13'b1101100011011,
13'b1101100011100,
13'b1101100101010,
13'b1101100101011,
13'b1101100101100,
13'b1101100101101,
13'b1101100111010,
13'b1101100111011,
13'b1101100111100,
13'b1110011011010,
13'b1110011011011,
13'b1110011101010,
13'b1110011101011,
13'b1110011101100,
13'b1110011111010,
13'b1110011111011,
13'b1110011111100,
13'b1110100001010,
13'b1110100001011,
13'b1110100001100,
13'b1110100001101,
13'b1110100011010,
13'b1110100011011,
13'b1110100011100,
13'b1110100011101,
13'b1110100101011,
13'b1110100101100,
13'b1110100101101,
13'b1110100111011,
13'b1110100111100,
13'b1110100111101,
13'b1111011101011,
13'b1111011101100,
13'b1111011111011,
13'b1111011111100,
13'b1111011111101,
13'b1111100001011,
13'b1111100001100,
13'b1111100001101,
13'b1111100011011,
13'b1111100011100,
13'b1111100011101,
13'b1111100101011,
13'b1111100101100,
13'b1111100101101,
13'b1111100111100,
13'b1111100111101: edge_mask_reg_512p3[86] <= 1'b1;
 		default: edge_mask_reg_512p3[86] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010100,
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100100,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110100,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000100,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010100,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100100,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100100,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110100,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000100,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010100,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100100,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1010010100,
13'b1010010101,
13'b1010010110,
13'b1010100100,
13'b1010100101,
13'b1010100110,
13'b1010110100,
13'b1010110101,
13'b1010110110,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b101010100100,
13'b101010100101,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b110010110100,
13'b110010110101,
13'b110011000100,
13'b110011000101,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b1000011010000,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1011011010000,
13'b1011011010001,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100100000,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1100011100000,
13'b1100011100001,
13'b1100011110000,
13'b1100011110001,
13'b1100100000000,
13'b1100100000001,
13'b1100100000010,
13'b1100100010000,
13'b1100100010001,
13'b1100100010010,
13'b1100100100000,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1101100000000,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100100000,
13'b1101100100001,
13'b1101100100010,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1110100010000,
13'b1110100100000,
13'b1110100110000,
13'b1110100110001,
13'b1110101000000,
13'b1110101000001,
13'b1110101000010,
13'b1110101010000,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101100000,
13'b1110101100010,
13'b1111100110000,
13'b1111101000000,
13'b1111101000001,
13'b1111101010000,
13'b1111101010001: edge_mask_reg_512p3[87] <= 1'b1;
 		default: edge_mask_reg_512p3[87] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011110101,
13'b10011110110,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b101100000101,
13'b101100000110,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111010101,
13'b110111010110,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101100000,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1100101110000,
13'b1100101110001,
13'b1100101110010,
13'b1100101110011,
13'b1100110000000,
13'b1100110000001,
13'b1100110000010,
13'b1100110000011,
13'b1100110010000,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110100000,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1101101110000,
13'b1101101110001,
13'b1101101110010,
13'b1101101110011,
13'b1101110000000,
13'b1101110000001,
13'b1101110000010,
13'b1101110000011,
13'b1101110010000,
13'b1101110010001,
13'b1101110010010,
13'b1101110010011,
13'b1101110100000,
13'b1101110100001,
13'b1101110100010,
13'b1101110100011,
13'b1101110110001,
13'b1101110110010,
13'b1101110110011,
13'b1110101000000,
13'b1110101000001,
13'b1110101000010,
13'b1110101010000,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101100000,
13'b1110101100001,
13'b1110101100010,
13'b1110101110000,
13'b1110101110001,
13'b1110101110010,
13'b1110110000000,
13'b1110110000001,
13'b1110110000010,
13'b1110110010000,
13'b1110110010001,
13'b1110110010010,
13'b1110110100000,
13'b1110110100001,
13'b1110110100010,
13'b1111101000000,
13'b1111101000001,
13'b1111101010000,
13'b1111101010001,
13'b1111101100000,
13'b1111101100001,
13'b1111101110000,
13'b1111101110001,
13'b1111110000000,
13'b1111110000001,
13'b1111110010000,
13'b1111110010001,
13'b1111110100000,
13'b1111110100001: edge_mask_reg_512p3[88] <= 1'b1;
 		default: edge_mask_reg_512p3[88] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11000101,
13'b11010100,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100100,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010100,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100100,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b100011100100,
13'b100011100101,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b110100000100,
13'b110100000101,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100100000,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1100100010000,
13'b1100100010001,
13'b1100100100000,
13'b1100100100001,
13'b1100100100010,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1101100100000,
13'b1101100100001,
13'b1101100100010,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1110100110000,
13'b1110100110001,
13'b1110101000000,
13'b1110101000001,
13'b1110101000010,
13'b1110101010000,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101100000,
13'b1110101100010,
13'b1111101000000,
13'b1111101000001,
13'b1111101010000,
13'b1111101010001: edge_mask_reg_512p3[89] <= 1'b1;
 		default: edge_mask_reg_512p3[89] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011110101,
13'b10011110110,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110101,
13'b11110110110,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110101,
13'b100110110110,
13'b101100000101,
13'b101100000110,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110101,
13'b101110110110,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110010101,
13'b110110010110,
13'b110110100101,
13'b110110100110,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000010,
13'b1000110000011,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101100000,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101100000,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1100101110000,
13'b1100101110001,
13'b1100101110010,
13'b1100101110011,
13'b1100110000001,
13'b1100110000010,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1101101110000,
13'b1101101110001,
13'b1101101110010,
13'b1101101110011,
13'b1101110000010,
13'b1110101000000,
13'b1110101000001,
13'b1110101000010,
13'b1110101010000,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101100000,
13'b1110101100001,
13'b1110101100010,
13'b1111101000000,
13'b1111101000001,
13'b1111101010000,
13'b1111101010001,
13'b1111101100000: edge_mask_reg_512p3[90] <= 1'b1;
 		default: edge_mask_reg_512p3[90] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010100,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010011,
13'b11100010100,
13'b11100010110,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110100100,
13'b11110100101,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110100100,
13'b100110100101,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101100000,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101100000,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1110101000000,
13'b1110101000001,
13'b1110101000010,
13'b1110101010000,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101100000,
13'b1110101100010,
13'b1111101000000,
13'b1111101000001,
13'b1111101010000,
13'b1111101010001: edge_mask_reg_512p3[91] <= 1'b1;
 		default: edge_mask_reg_512p3[91] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1010100101,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b11010110101,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b100010110101,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b111011100100,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b1000011100011,
13'b1000011100100,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1001011100010,
13'b1001011100011,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1011011100010,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100100000,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1100011100001,
13'b1100011100010,
13'b1100011110000,
13'b1100011110001,
13'b1100011110010,
13'b1100100000000,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100010000,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100100000,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1101011110001,
13'b1101011110010,
13'b1101100000000,
13'b1101100000001,
13'b1101100000010,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100100000,
13'b1101100100001,
13'b1101100100010,
13'b1101100100011,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1110100000000,
13'b1110100000001,
13'b1110100010000,
13'b1110100010001,
13'b1110100100000,
13'b1110100100001,
13'b1110100110000,
13'b1110100110001,
13'b1110100110010,
13'b1110101000000,
13'b1110101000001,
13'b1110101000010,
13'b1110101010000,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101100000,
13'b1110101100010,
13'b1111100100000,
13'b1111100110000,
13'b1111101000000,
13'b1111101000001,
13'b1111101010000,
13'b1111101010001: edge_mask_reg_512p3[92] <= 1'b1;
 		default: edge_mask_reg_512p3[92] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[93] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[94] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000110100101,
13'b1000110100110,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110001,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1011110100100,
13'b1011110100101,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111110001,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1100110100100,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111110001,
13'b1100111110010,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1101111010001,
13'b1101111010010,
13'b1101111010011,
13'b1101111100001,
13'b1101111100010,
13'b1101111100011,
13'b1101111100100,
13'b1101111110001,
13'b1101111110010,
13'b1101111110011,
13'b1101111110100: edge_mask_reg_512p3[95] <= 1'b1;
 		default: edge_mask_reg_512p3[95] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100100101001,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101011000,
13'b110101011001,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101110111,
13'b1000101111000,
13'b1000101111001,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1000110010111,
13'b1000110011000,
13'b1000110011001,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111001001,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110111,
13'b1001101111000,
13'b1001101111001,
13'b1001110000111,
13'b1001110001000,
13'b1001110001001,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110011001,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110101001,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001110111001,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010101011000,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110111,
13'b1010101111000,
13'b1010101111001,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110001001,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1010110011001,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010110111000,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111011000,
13'b1010111100110,
13'b1010111100111,
13'b1010111101000,
13'b1011101011000,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011110111000,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111001000,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111011000,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110101,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1100110010100,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1100110100100,
13'b1100110100101,
13'b1100110100110,
13'b1100110100111,
13'b1100110101000,
13'b1100110110100,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100110111000,
13'b1100111000100,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111001000,
13'b1100111010100,
13'b1100111010101,
13'b1100111010110,
13'b1100111010111,
13'b1100111100101,
13'b1100111100110,
13'b1100111100111,
13'b1101101100101,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110100,
13'b1101101110101,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101110000100,
13'b1101110000101,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1101110010100,
13'b1101110010101,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1101110100111,
13'b1101110101000,
13'b1101110110100,
13'b1101110110101,
13'b1101110110110,
13'b1101110110111,
13'b1101110111000,
13'b1101111000100,
13'b1101111000101,
13'b1101111000110,
13'b1101111000111,
13'b1101111010100,
13'b1101111010101,
13'b1101111010110,
13'b1101111010111,
13'b1101111100110,
13'b1101111100111,
13'b1110101100101,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110100,
13'b1110101110101,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110110000100,
13'b1110110000101,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110010100,
13'b1110110010101,
13'b1110110010110,
13'b1110110010111,
13'b1110110011000,
13'b1110110100100,
13'b1110110100101,
13'b1110110100110,
13'b1110110100111,
13'b1110110110100,
13'b1110110110101,
13'b1110110110111,
13'b1110111000100,
13'b1111101110101,
13'b1111101110110,
13'b1111110000101,
13'b1111110000110,
13'b1111110010100,
13'b1111110010101: edge_mask_reg_512p3[96] <= 1'b1;
 		default: edge_mask_reg_512p3[96] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b100000110000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000110,
13'b100001000111,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000110,
13'b101001000111,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000110,
13'b110001000111,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010110,
13'b111000100000,
13'b111000100001: edge_mask_reg_512p3[97] <= 1'b1;
 		default: edge_mask_reg_512p3[97] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[98] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011110101,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b101100000101,
13'b101100000110,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111010101,
13'b110111010110,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1011100110000,
13'b1011100110001,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101100000,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1100101000000,
13'b1100101010000,
13'b1100101010001,
13'b1100101100000,
13'b1100101100001,
13'b1100101100010,
13'b1100101110000,
13'b1100101110001,
13'b1100101110010,
13'b1100110000000,
13'b1100110000001,
13'b1100110000010,
13'b1100110000011,
13'b1100110010000,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110100000,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1101101010000,
13'b1101101100000,
13'b1101101100001,
13'b1101101110000,
13'b1101101110001,
13'b1101101110010,
13'b1101110000000,
13'b1101110000001,
13'b1101110000010,
13'b1101110010000,
13'b1101110010001,
13'b1101110010010,
13'b1101110010011,
13'b1101110100000,
13'b1101110100001,
13'b1101110100010,
13'b1101110100011,
13'b1101110110001,
13'b1101110110010,
13'b1101110110011,
13'b1110101100000,
13'b1110101110000,
13'b1110101110001,
13'b1110110000000,
13'b1110110000001,
13'b1110110010000,
13'b1110110010001,
13'b1110110010010,
13'b1110110100000,
13'b1110110100001,
13'b1110110100010,
13'b1111101110000,
13'b1111110000000,
13'b1111110010000,
13'b1111110010001,
13'b1111110100000,
13'b1111110100001: edge_mask_reg_512p3[99] <= 1'b1;
 		default: edge_mask_reg_512p3[99] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011110101,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101100000101,
13'b101100000110,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010101,
13'b101111010110,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000101,
13'b110111000110,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100011,
13'b1000110100100,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110100010,
13'b1001110100011,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1011100110000,
13'b1011100110001,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101100000,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110100010,
13'b1011110100011,
13'b1100101000000,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101100000,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1100101110000,
13'b1100101110001,
13'b1100101110010,
13'b1100101110011,
13'b1100110000000,
13'b1100110000001,
13'b1100110000010,
13'b1100110000011,
13'b1100110010000,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110100010,
13'b1100110100011,
13'b1101101010000,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1101101110000,
13'b1101101110001,
13'b1101101110010,
13'b1101101110011,
13'b1101110000000,
13'b1101110000001,
13'b1101110000010,
13'b1101110000011,
13'b1101110010000,
13'b1101110010001,
13'b1101110010010,
13'b1101110010011,
13'b1101110100010,
13'b1110101010000,
13'b1110101100000,
13'b1110101100001,
13'b1110101110000,
13'b1110101110001,
13'b1110110000000,
13'b1110110000001,
13'b1110110000010,
13'b1110110010000,
13'b1110110010001,
13'b1110110010010,
13'b1111101100000,
13'b1111101110000,
13'b1111101110001,
13'b1111110000000,
13'b1111110000001,
13'b1111110010000,
13'b1111110010001: edge_mask_reg_512p3[100] <= 1'b1;
 		default: edge_mask_reg_512p3[100] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b100011111000,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110001000,
13'b110110001001,
13'b111100100111,
13'b111100101000,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101111000,
13'b111101111001,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101110111,
13'b1000101111000,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110111,
13'b1001101111000,
13'b1010100100111,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110111,
13'b1010101111000,
13'b1011100100110,
13'b1011100100111,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110111,
13'b1011101111000,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110111,
13'b1100101111000,
13'b1101100100111,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110110,
13'b1101101110111,
13'b1110100110101,
13'b1110100110110,
13'b1110100110111,
13'b1110101000101,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101010101,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110111,
13'b1111100110101,
13'b1111100110110,
13'b1111100110111,
13'b1111101000101,
13'b1111101000110,
13'b1111101000111,
13'b1111101001000,
13'b1111101010101,
13'b1111101010110,
13'b1111101010111,
13'b1111101011000,
13'b1111101100110,
13'b1111101100111: edge_mask_reg_512p3[101] <= 1'b1;
 		default: edge_mask_reg_512p3[101] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[102] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100101101001,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110010111,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000110010111,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110010111,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010110010110,
13'b1010110010111,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010110111000,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111011000,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111101000,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1010111111000,
13'b1011110010110,
13'b1011110010111,
13'b1011110100101,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110101,
13'b1011111110110,
13'b1011111110111,
13'b1100110100101,
13'b1100110100110,
13'b1100110100111,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111010101,
13'b1100111010110,
13'b1100111010111,
13'b1100111100101,
13'b1100111100110,
13'b1100111100111,
13'b1100111110101,
13'b1100111110110,
13'b1100111110111,
13'b1101110100101,
13'b1101110100110,
13'b1101110100111,
13'b1101110110101,
13'b1101110110110,
13'b1101110110111,
13'b1101111000101,
13'b1101111000110,
13'b1101111000111,
13'b1101111010101,
13'b1101111010110,
13'b1101111010111,
13'b1101111100101,
13'b1101111100110,
13'b1101111100111,
13'b1101111110101,
13'b1101111110110,
13'b1101111110111,
13'b1110110100101,
13'b1110110100110,
13'b1110110110101,
13'b1110110110110,
13'b1110110110111,
13'b1110111000101,
13'b1110111000110,
13'b1110111000111,
13'b1110111010101,
13'b1110111010110,
13'b1110111100100,
13'b1110111100101,
13'b1110111100110,
13'b1110111110100,
13'b1110111110101,
13'b1110111110110,
13'b1111110100101,
13'b1111110110101,
13'b1111110110110,
13'b1111111000101,
13'b1111111000110,
13'b1111111010100,
13'b1111111010101,
13'b1111111010110,
13'b1111111100100,
13'b1111111100101,
13'b1111111100110,
13'b1111111110100,
13'b1111111110101,
13'b1111111110110: edge_mask_reg_512p3[103] <= 1'b1;
 		default: edge_mask_reg_512p3[103] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100101011010,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b101111011011,
13'b110110000111,
13'b110110001000,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110000111,
13'b111110001000,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001110111001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010110000110,
13'b1010110000111,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010110111000,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110010,
13'b1010111110100,
13'b1010111110101,
13'b1011110000110,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011110111000,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1100110100100,
13'b1100110100101,
13'b1100110100110,
13'b1100110100111,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111010011,
13'b1100111010100,
13'b1100111100011,
13'b1101110010101,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1101110110011,
13'b1101110110100,
13'b1101110110101,
13'b1101110110110,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111010011,
13'b1101111010100,
13'b1110110100100,
13'b1110110100101,
13'b1110110110100,
13'b1110110110101,
13'b1110111000100: edge_mask_reg_512p3[104] <= 1'b1;
 		default: edge_mask_reg_512p3[104] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100111000,
13'b100111001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b11001001001,
13'b11001001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b100001001001,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110101,
13'b101001110110,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011111000,
13'b110011111001,
13'b110100001000,
13'b110100001001,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1001001110100,
13'b1001001110101,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011100010,
13'b1010011100011,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010110010,
13'b1011010110011,
13'b1011010110100,
13'b1011011000010,
13'b1011011000011,
13'b1011011010010,
13'b1011011010011,
13'b1011011100010,
13'b1100010000011,
13'b1100010010011,
13'b1100010100011,
13'b1100010110011,
13'b1100011000011,
13'b1100011010011: edge_mask_reg_512p3[105] <= 1'b1;
 		default: edge_mask_reg_512p3[105] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b10001111001,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010011000,
13'b110010011001,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010101000,
13'b110010101001,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1001010110010,
13'b1001010110011,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100100,
13'b1001100100101,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1011011000010,
13'b1011011000011,
13'b1011011010010,
13'b1011011010011,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010011,
13'b1011100010100,
13'b1100011010011,
13'b1100011100011,
13'b1100011110011,
13'b1100011110100,
13'b1100100000011,
13'b1100100000100,
13'b1100100010011,
13'b1100100010100: edge_mask_reg_512p3[106] <= 1'b1;
 		default: edge_mask_reg_512p3[106] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100100111001,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b101111011011,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101111000,
13'b111101111001,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110101000,
13'b111110101001,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000101111000,
13'b1000101111001,
13'b1000110001000,
13'b1000110001001,
13'b1000110010111,
13'b1000110011000,
13'b1000110011001,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000111000111,
13'b1000111001000,
13'b1000111001001,
13'b1000111010111,
13'b1000111011000,
13'b1000111011001,
13'b1000111100111,
13'b1000111101000,
13'b1000111101001,
13'b1001101111000,
13'b1001101111001,
13'b1001110000111,
13'b1001110001000,
13'b1001110001001,
13'b1001110010111,
13'b1001110011000,
13'b1001110011001,
13'b1001110100111,
13'b1001110101000,
13'b1001110101001,
13'b1001110110111,
13'b1001110111000,
13'b1001110111001,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111001001,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111011001,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010101110111,
13'b1010101111000,
13'b1010101111001,
13'b1010110000111,
13'b1010110001000,
13'b1010110001001,
13'b1010110010111,
13'b1010110011000,
13'b1010110011001,
13'b1010110100111,
13'b1010110101000,
13'b1010110101001,
13'b1010110110110,
13'b1010110110111,
13'b1010110111000,
13'b1010110111001,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111001001,
13'b1010111010110,
13'b1010111010111,
13'b1010111011000,
13'b1010111100110,
13'b1010111100111,
13'b1010111101000,
13'b1010111110111,
13'b1011101110111,
13'b1011101111000,
13'b1011101111001,
13'b1011110000111,
13'b1011110001000,
13'b1011110001001,
13'b1011110010111,
13'b1011110011000,
13'b1011110011001,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110101001,
13'b1011110110110,
13'b1011110110111,
13'b1011110111000,
13'b1011110111001,
13'b1011111000110,
13'b1011111000111,
13'b1011111001000,
13'b1011111010110,
13'b1011111010111,
13'b1011111011000,
13'b1011111100110,
13'b1011111100111,
13'b1011111101000,
13'b1011111110111,
13'b1100101110111,
13'b1100101111000,
13'b1100101111001,
13'b1100110000111,
13'b1100110001000,
13'b1100110001001,
13'b1100110010111,
13'b1100110011000,
13'b1100110011001,
13'b1100110100110,
13'b1100110100111,
13'b1100110101000,
13'b1100110101001,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100110111000,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111001000,
13'b1100111010101,
13'b1100111010110,
13'b1100111010111,
13'b1100111011000,
13'b1100111100110,
13'b1100111100111,
13'b1100111101000,
13'b1100111110111,
13'b1101101110111,
13'b1101101111000,
13'b1101101111001,
13'b1101110000111,
13'b1101110001000,
13'b1101110001001,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1101110011001,
13'b1101110100110,
13'b1101110100111,
13'b1101110101000,
13'b1101110101001,
13'b1101110110101,
13'b1101110110110,
13'b1101110110111,
13'b1101110111000,
13'b1101111000101,
13'b1101111000110,
13'b1101111000111,
13'b1101111001000,
13'b1101111010101,
13'b1101111010110,
13'b1101111010111,
13'b1101111011000,
13'b1101111100110,
13'b1101111100111,
13'b1110101110111,
13'b1110101111000,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110010110,
13'b1110110010111,
13'b1110110011000,
13'b1110110100101,
13'b1110110100110,
13'b1110110100111,
13'b1110110101000,
13'b1110110110101,
13'b1110110110110,
13'b1110110110111,
13'b1110110111000,
13'b1110111000101,
13'b1110111000110,
13'b1110111000111,
13'b1110111010101,
13'b1110111010110,
13'b1110111010111,
13'b1111110000110,
13'b1111110000111,
13'b1111110001000,
13'b1111110010110,
13'b1111110010111,
13'b1111110011000,
13'b1111110100101,
13'b1111110100110,
13'b1111110100111,
13'b1111110101000,
13'b1111110110101,
13'b1111110110110,
13'b1111110110111,
13'b1111111000101,
13'b1111111000110,
13'b1111111000111,
13'b1111111010101,
13'b1111111010110: edge_mask_reg_512p3[107] <= 1'b1;
 		default: edge_mask_reg_512p3[107] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100101000101,
13'b100101000110,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101101000110,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111110001,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111010000,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111110001,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1100110000000,
13'b1100110010000,
13'b1100110010001,
13'b1100110100000,
13'b1100110100001,
13'b1100110100010,
13'b1100110110000,
13'b1100110110001,
13'b1100110110010,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111010000,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111100000,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111110001,
13'b1100111110010,
13'b1100111110011,
13'b1101110010000,
13'b1101110100000,
13'b1101110100001,
13'b1101110110000,
13'b1101110110001,
13'b1101111000000,
13'b1101111000001,
13'b1101111000010,
13'b1101111010000,
13'b1101111010001,
13'b1101111010010,
13'b1101111100000,
13'b1101111100001,
13'b1101111100010,
13'b1101111100011,
13'b1101111110000,
13'b1101111110001,
13'b1101111110010,
13'b1101111110011,
13'b1110110100000,
13'b1110110110000,
13'b1110110110001,
13'b1110111000000,
13'b1110111000001,
13'b1110111010000,
13'b1110111010001,
13'b1110111010010,
13'b1110111100000,
13'b1110111100001,
13'b1110111100010,
13'b1110111110000,
13'b1110111110001,
13'b1110111110010,
13'b1111111000001,
13'b1111111010001,
13'b1111111010010,
13'b1111111100001,
13'b1111111100010,
13'b1111111110001,
13'b1111111110010: edge_mask_reg_512p3[108] <= 1'b1;
 		default: edge_mask_reg_512p3[108] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[109] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110101110110,
13'b110101110111,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110000,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1010110010001,
13'b1010110010010,
13'b1010110100001,
13'b1010110100010,
13'b1010110110001,
13'b1010110110010,
13'b1010111000001,
13'b1010111000010,
13'b1010111010001,
13'b1010111010010,
13'b1010111100001,
13'b1010111100010,
13'b1010111110001,
13'b1010111110010: edge_mask_reg_512p3[110] <= 1'b1;
 		default: edge_mask_reg_512p3[110] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10110000110,
13'b10110000111,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110010,
13'b11110110011,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100010,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110110010110,
13'b110110010111,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111110110000,
13'b111110110001,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000110,
13'b111111000111,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010110,
13'b111111010111,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100110,
13'b111111100111,
13'b1000111010000,
13'b1000111010001,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011: edge_mask_reg_512p3[111] <= 1'b1;
 		default: edge_mask_reg_512p3[111] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111000110,
13'b100111000111,
13'b101111000110,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111111100010: edge_mask_reg_512p3[112] <= 1'b1;
 		default: edge_mask_reg_512p3[112] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101101000,
13'b101101001,
13'b101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101111010,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100110001010,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101110101001,
13'b101110101010,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110111001,
13'b101110111010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b101111011011,
13'b110111000100,
13'b110111000101,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b111111100011,
13'b111111100100,
13'b111111100101: edge_mask_reg_512p3[113] <= 1'b1;
 		default: edge_mask_reg_512p3[113] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b1001101001,
13'b1001101010,
13'b1001111001,
13'b1001111010,
13'b1010001001,
13'b1010001010,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100000,
13'b11001100001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110000,
13'b11001110001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000000,
13'b11010000001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100000,
13'b100001100001,
13'b100001100010,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110000,
13'b100001110001,
13'b100001110010,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000000,
13'b100010000001,
13'b100010000010,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010000,
13'b100010010001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b101000100111,
13'b101000101000,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100000,
13'b101010100001,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b110000110111,
13'b110000111000,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100001,
13'b110010100100,
13'b110010100101,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b111001000011,
13'b111001000100,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1001001010010,
13'b1001001010011,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100010,
13'b1001010100011,
13'b1010001100011,
13'b1010001110010,
13'b1010001110011,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100: edge_mask_reg_512p3[114] <= 1'b1;
 		default: edge_mask_reg_512p3[114] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001101010,
13'b10001101011,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001101010,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001011010,
13'b101000101001,
13'b101000101010,
13'b101000101011,
13'b101000111001,
13'b101000111010,
13'b111000011001,
13'b111000011010,
13'b111000011011,
13'b111000011100,
13'b111000101010,
13'b111000101011,
13'b1000000011001,
13'b1000000011010,
13'b1000000011011,
13'b1000000011100,
13'b1000000101010,
13'b1000000101011,
13'b1000000101100,
13'b1001000011001,
13'b1001000011010,
13'b1001000011011,
13'b1001000011100,
13'b1001000101011,
13'b1001000101100,
13'b1010000001001,
13'b1010000001010,
13'b1010000001011,
13'b1010000001100,
13'b1010000011001,
13'b1010000011010,
13'b1010000011011,
13'b1010000011100,
13'b1010000101011,
13'b1010000101100,
13'b1011000001001,
13'b1011000001010,
13'b1011000001011,
13'b1011000001100,
13'b1011000011001,
13'b1011000011010,
13'b1011000011011,
13'b1011000011100,
13'b1011000101010,
13'b1011000101011,
13'b1011000101100,
13'b1100000001001,
13'b1100000001010,
13'b1100000001011,
13'b1100000001100,
13'b1100000011001,
13'b1100000011010,
13'b1100000011011,
13'b1100000011100,
13'b1100000101010,
13'b1100000101011,
13'b1100000101100,
13'b1101000001001,
13'b1101000001010,
13'b1101000001011,
13'b1101000001100,
13'b1101000011001,
13'b1101000011010,
13'b1101000011011,
13'b1101000011100,
13'b1101000101011,
13'b1101000101100,
13'b1110000001001,
13'b1110000001010,
13'b1110000001011,
13'b1110000001100,
13'b1110000011010,
13'b1110000011011,
13'b1110000011100,
13'b1111000001001,
13'b1111000001010,
13'b1111000001011,
13'b1111000001100,
13'b1111000011010,
13'b1111000011011,
13'b1111000011100: edge_mask_reg_512p3[115] <= 1'b1;
 		default: edge_mask_reg_512p3[115] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100010110,
13'b1100010111,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100100100110,
13'b100100100111,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100100111,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000010,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000101010001,
13'b1000101010010,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1001101100001,
13'b1001101100010,
13'b1001101110001,
13'b1001101110010,
13'b1001110000001,
13'b1001110000010,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1010110110001,
13'b1010110110010,
13'b1010111000001,
13'b1010111000010,
13'b1010111010001,
13'b1010111010010,
13'b1010111100001,
13'b1010111100010: edge_mask_reg_512p3[116] <= 1'b1;
 		default: edge_mask_reg_512p3[116] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101110111,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101110111,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111100000,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1011110100010,
13'b1011110100011,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111010000,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111100000,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111010000,
13'b1100111010010,
13'b1100111010011: edge_mask_reg_512p3[117] <= 1'b1;
 		default: edge_mask_reg_512p3[117] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000111000,
13'b100000111001,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b1010000000011,
13'b1010000000100: edge_mask_reg_512p3[118] <= 1'b1;
 		default: edge_mask_reg_512p3[118] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[119] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[120] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[121] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101110000111,
13'b101110001000,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110110110,
13'b1000110110111,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001110110110,
13'b1001110110111,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110001,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1011111100000,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111110000,
13'b1011111110001,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1100110110100,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111010000,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111010110,
13'b1100111010111,
13'b1100111100000,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111100110,
13'b1100111110000,
13'b1100111110001,
13'b1100111110010,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1101110110011,
13'b1101110110100,
13'b1101110110101,
13'b1101110110110,
13'b1101111000001,
13'b1101111000010,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111000110,
13'b1101111000111,
13'b1101111010000,
13'b1101111010001,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1101111010101,
13'b1101111010110,
13'b1101111100000,
13'b1101111100001,
13'b1101111100010,
13'b1101111100011,
13'b1101111100100,
13'b1101111100101,
13'b1101111100110,
13'b1101111110000,
13'b1101111110001,
13'b1101111110010,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1110110110010,
13'b1110110110011,
13'b1110110110100,
13'b1110110110101,
13'b1110110110110,
13'b1110111000001,
13'b1110111000010,
13'b1110111000011,
13'b1110111000100,
13'b1110111000101,
13'b1110111000110,
13'b1110111000111,
13'b1110111010001,
13'b1110111010010,
13'b1110111010011,
13'b1110111010100,
13'b1110111010101,
13'b1110111010110,
13'b1110111100000,
13'b1110111100001,
13'b1110111100010,
13'b1110111100011,
13'b1110111100100,
13'b1110111100101,
13'b1110111110000,
13'b1110111110001,
13'b1110111110010,
13'b1111110110011,
13'b1111110110100,
13'b1111110110101,
13'b1111111000010,
13'b1111111000011,
13'b1111111000100,
13'b1111111000101,
13'b1111111010001,
13'b1111111010010,
13'b1111111010011,
13'b1111111010100,
13'b1111111010101,
13'b1111111100001,
13'b1111111100010: edge_mask_reg_512p3[122] <= 1'b1;
 		default: edge_mask_reg_512p3[122] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100110101010,
13'b100110101011,
13'b100110110110,
13'b100110111010,
13'b100110111011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110111000101,
13'b110111010100,
13'b110111010101,
13'b110111010110: edge_mask_reg_512p3[123] <= 1'b1;
 		default: edge_mask_reg_512p3[123] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1001111001,
13'b1001111010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101100100,
13'b10101100101,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011010,
13'b10110011011,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100100,
13'b100101100101,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001010,
13'b101010101001,
13'b101010101010,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101100100,
13'b101101100101,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011010,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101010,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100110010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010010,
13'b1000100010011,
13'b1001011000010,
13'b1001011000011,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001100000010,
13'b1001100000011,
13'b1010011010010,
13'b1010011010011,
13'b1010011100010,
13'b1010011100011,
13'b1010011110011: edge_mask_reg_512p3[124] <= 1'b1;
 		default: edge_mask_reg_512p3[124] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011001,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101001001,
13'b110101010011,
13'b110101010100,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110011000,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110101000,
13'b111110101001,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110111000,
13'b111110111001,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111001000,
13'b111111001001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b1000110100000,
13'b1000110110000,
13'b1000110110001: edge_mask_reg_512p3[125] <= 1'b1;
 		default: edge_mask_reg_512p3[125] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100011001000,
13'b100011001001,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000000,
13'b100100000001,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010000,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100000,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000000,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010000,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110011011000,
13'b110011011001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011101000,
13'b110011101001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111000,
13'b110011111001,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101111001,
13'b110101111010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b111011110010,
13'b111011110011,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100001000,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100011000,
13'b111100011001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100101000,
13'b111100101001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010011,
13'b111101010100,
13'b111101100011,
13'b111101100100,
13'b111101110011,
13'b111101110100,
13'b1000100100011,
13'b1000100110011: edge_mask_reg_512p3[126] <= 1'b1;
 		default: edge_mask_reg_512p3[126] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110001,
13'b11110010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000001,
13'b100000010,
13'b100000011,
13'b100000100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010001,
13'b100010010,
13'b100010011,
13'b100010100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100001,
13'b100100010,
13'b100100011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110001,
13'b100110010,
13'b100110011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000001,
13'b101000010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010011,
13'b1011010100,
13'b1011010101,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100011,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110001,
13'b1011110010,
13'b1011110011,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000001,
13'b1100000010,
13'b1100000011,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010001,
13'b1100010010,
13'b1100010011,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100001,
13'b1100100010,
13'b1100100011,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110001,
13'b1100110010,
13'b1100110011,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000001,
13'b1101000010,
13'b1101000011,
13'b1101000100,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010001,
13'b1101010010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10010111001,
13'b10010111010,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010001,
13'b10100010010,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100001,
13'b10100100010,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110001,
13'b10100110010,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000001,
13'b10101000010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010001,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100001,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110100001001,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010,
13'b110100111001,
13'b110100111010,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101011001,
13'b110101011010,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101101001,
13'b110101101010,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101111001,
13'b110101111010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110: edge_mask_reg_512p3[127] <= 1'b1;
 		default: edge_mask_reg_512p3[127] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101010,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b111101001001,
13'b111101001010,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110001001,
13'b111110001010,
13'b1000101001001,
13'b1000101001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101011010,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1000110001001,
13'b1000110001010,
13'b1000110001011,
13'b1001101001001,
13'b1001101001010,
13'b1001101011000,
13'b1001101011001,
13'b1001101011010,
13'b1001101101001,
13'b1001101101010,
13'b1001101101011,
13'b1001101111001,
13'b1001101111010,
13'b1001101111011,
13'b1001110001001,
13'b1001110001010,
13'b1001110001011,
13'b1010101001000,
13'b1010101001001,
13'b1010101001010,
13'b1010101011000,
13'b1010101011001,
13'b1010101011010,
13'b1010101101000,
13'b1010101101001,
13'b1010101101010,
13'b1010101101011,
13'b1010101111000,
13'b1010101111001,
13'b1010101111010,
13'b1010101111011,
13'b1010110001001,
13'b1010110001010,
13'b1010110001011,
13'b1011101001000,
13'b1011101001001,
13'b1011101001010,
13'b1011101011000,
13'b1011101011001,
13'b1011101011010,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1011101101010,
13'b1011101110111,
13'b1011101111000,
13'b1011101111001,
13'b1011101111010,
13'b1011101111011,
13'b1011110001001,
13'b1011110001010,
13'b1100101001000,
13'b1100101001001,
13'b1100101001010,
13'b1100101011000,
13'b1100101011001,
13'b1100101011010,
13'b1100101100111,
13'b1100101101000,
13'b1100101101001,
13'b1100101101010,
13'b1100101101011,
13'b1100101110111,
13'b1100101111000,
13'b1100101111001,
13'b1100101111010,
13'b1100101111011,
13'b1100110000111,
13'b1100110001000,
13'b1100110001001,
13'b1100110001010,
13'b1100110001011,
13'b1101101001001,
13'b1101101011000,
13'b1101101011001,
13'b1101101011010,
13'b1101101100111,
13'b1101101101000,
13'b1101101101001,
13'b1101101101010,
13'b1101101110111,
13'b1101101111000,
13'b1101101111001,
13'b1101101111010,
13'b1101110000111,
13'b1101110001000,
13'b1101110001001,
13'b1101110001010,
13'b1110101100111,
13'b1110101101000,
13'b1110101101001,
13'b1110101101010,
13'b1110101110111,
13'b1110101111000,
13'b1110101111001,
13'b1110101111010,
13'b1110110000111,
13'b1110110001000,
13'b1110110001001,
13'b1111101100111,
13'b1111101101000,
13'b1111101101001,
13'b1111101110111,
13'b1111101111000,
13'b1111101111001,
13'b1111110000111,
13'b1111110001000: edge_mask_reg_512p3[128] <= 1'b1;
 		default: edge_mask_reg_512p3[128] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100111001,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b1000101111000,
13'b1000101111001,
13'b1000101111010,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1000110001010,
13'b1000110010111,
13'b1000110011000,
13'b1000110011001,
13'b1000110011010,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110101010,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000111000111,
13'b1000111001000,
13'b1001101111000,
13'b1001101111001,
13'b1001101111010,
13'b1001110000111,
13'b1001110001000,
13'b1001110001001,
13'b1001110001010,
13'b1001110010111,
13'b1001110011000,
13'b1001110011001,
13'b1001110011010,
13'b1001110100111,
13'b1001110101000,
13'b1001110101001,
13'b1001110101010,
13'b1001110110111,
13'b1001110111000,
13'b1001110111001,
13'b1001111000111,
13'b1001111001000,
13'b1001111001001,
13'b1010101111000,
13'b1010101111001,
13'b1010101111010,
13'b1010110000111,
13'b1010110001000,
13'b1010110001001,
13'b1010110001010,
13'b1010110010111,
13'b1010110011000,
13'b1010110011001,
13'b1010110011010,
13'b1010110100111,
13'b1010110101000,
13'b1010110101001,
13'b1010110101010,
13'b1010110110111,
13'b1010110111000,
13'b1010110111001,
13'b1010111000111,
13'b1010111001000,
13'b1011101111000,
13'b1011101111001,
13'b1011101111010,
13'b1011110000111,
13'b1011110001000,
13'b1011110001001,
13'b1011110010111,
13'b1011110011000,
13'b1011110011001,
13'b1011110011010,
13'b1011110100111,
13'b1011110101000,
13'b1011110101001,
13'b1011110101010,
13'b1011110110111,
13'b1011110111000,
13'b1011110111001,
13'b1011111000111,
13'b1011111001000,
13'b1100101111000,
13'b1100101111001,
13'b1100101111010,
13'b1100110000111,
13'b1100110001000,
13'b1100110001001,
13'b1100110001010,
13'b1100110010111,
13'b1100110011000,
13'b1100110011001,
13'b1100110011010,
13'b1100110100111,
13'b1100110101000,
13'b1100110101001,
13'b1100110110111,
13'b1100110111000,
13'b1100110111001,
13'b1100111000111,
13'b1100111001000,
13'b1100111010111,
13'b1101101111000,
13'b1101101111001,
13'b1101101111010,
13'b1101110000111,
13'b1101110001000,
13'b1101110001001,
13'b1101110001010,
13'b1101110010111,
13'b1101110011000,
13'b1101110011001,
13'b1101110011010,
13'b1101110100110,
13'b1101110100111,
13'b1101110101000,
13'b1101110101001,
13'b1101110110110,
13'b1101110110111,
13'b1101110111000,
13'b1101110111001,
13'b1101111000110,
13'b1101111000111,
13'b1101111001000,
13'b1110101111000,
13'b1110101111001,
13'b1110101111010,
13'b1110110000111,
13'b1110110001000,
13'b1110110001001,
13'b1110110001010,
13'b1110110010111,
13'b1110110011000,
13'b1110110011001,
13'b1110110011010,
13'b1110110100110,
13'b1110110100111,
13'b1110110101000,
13'b1110110101001,
13'b1110110110110,
13'b1110110110111,
13'b1110110111000,
13'b1110110111001,
13'b1110111000110,
13'b1110111000111,
13'b1110111001000,
13'b1111101110111,
13'b1111101111000,
13'b1111101111001,
13'b1111110000111,
13'b1111110001000,
13'b1111110001001,
13'b1111110010110,
13'b1111110010111,
13'b1111110011000,
13'b1111110011001,
13'b1111110100110,
13'b1111110100111,
13'b1111110101000,
13'b1111110101001,
13'b1111110110110,
13'b1111110110111,
13'b1111110111000,
13'b1111110111001,
13'b1111111000111,
13'b1111111001000: edge_mask_reg_512p3[129] <= 1'b1;
 		default: edge_mask_reg_512p3[129] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[130] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110000,
13'b1011110111,
13'b1011111000,
13'b1100000111,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000000,
13'b10011000001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010000,
13'b10011010001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100000,
13'b10011100001,
13'b10011100010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110000,
13'b10011110001,
13'b10011110010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000000,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110100,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000000,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010000,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100000,
13'b11011100001,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110000,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000000,
13'b11100000001,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110001,
13'b100010110010,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110000,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000000,
13'b100100000001,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010000,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b101010100111,
13'b101010101000,
13'b101010110011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110000,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000000,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010000,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000100,
13'b101101000101,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b111011010010,
13'b111011010011,
13'b111011010111,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100111,
13'b111011101000,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b1000011100010,
13'b1000011100011,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000010,
13'b1000101000011,
13'b1001100000010,
13'b1001100000011,
13'b1001100010010,
13'b1001100010011,
13'b1001100100010,
13'b1001100100011,
13'b1001100110011: edge_mask_reg_512p3[131] <= 1'b1;
 		default: edge_mask_reg_512p3[131] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000111,
13'b1101001000,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000000,
13'b10011000001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010000,
13'b10011010001,
13'b10011010100,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100000,
13'b10011100001,
13'b10011100010,
13'b10011100100,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110000,
13'b10011110001,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100000,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110000,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000000,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010000,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100000,
13'b11011100001,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110000,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000000,
13'b11100000001,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b100000111000,
13'b100000111001,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000000,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010000,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100000,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110000,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000000,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110000,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000000,
13'b100100000001,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110111,
13'b100100111000,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000000,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110111,
13'b101100111000,
13'b110001001001,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001011000,
13'b110001011001,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001101000,
13'b110001101001,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000010,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010011000,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010101000,
13'b111010101001,
13'b111010110010,
13'b111010110011,
13'b111010111000,
13'b111010111001,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110111,
13'b111011111000,
13'b1000010000001: edge_mask_reg_512p3[132] <= 1'b1;
 		default: edge_mask_reg_512p3[132] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100111,
13'b1101110111,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10100000111,
13'b10100001000,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000000,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101100010111,
13'b101100011000,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010000,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100000,
13'b110110100100,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b111100110010,
13'b111100110011,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000111,
13'b111101001000,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110100000,
13'b111110100001,
13'b111110100011,
13'b111110100100,
13'b1000101000010,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100000,
13'b1000110100010,
13'b1000110100011,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100010,
13'b1010101110010,
13'b1010101110011,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010010,
13'b1010110010011: edge_mask_reg_512p3[133] <= 1'b1;
 		default: edge_mask_reg_512p3[133] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11010100111,
13'b11010101000,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b100010100111,
13'b100010101000,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100111,
13'b100110101000,
13'b101010101000,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000000,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011101000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011111000,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100001000,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100011001,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111110000010,
13'b111110000011,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101100010,
13'b1000101100011,
13'b1000101110010,
13'b1000101110011,
13'b1001011010010,
13'b1001011010011,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000010,
13'b1001101000011,
13'b1001101010010,
13'b1001101010011,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100110010,
13'b1010100110011,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011100000000,
13'b1011100000001: edge_mask_reg_512p3[134] <= 1'b1;
 		default: edge_mask_reg_512p3[134] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11010110,
13'b11010111,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101010110,
13'b1101010111,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10011100110,
13'b10011100111,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010000,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100000,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110000,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000000,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010000,
13'b11101010001,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100000,
13'b11101100001,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000010,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010000,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100000,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100111,
13'b100110101000,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000000,
13'b101100000001,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010000,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000000,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b110011110110,
13'b110011110111,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b111100100001,
13'b111100100110,
13'b111100100111,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b1000101100010,
13'b1000101100011,
13'b1000101110010,
13'b1000101110011: edge_mask_reg_512p3[135] <= 1'b1;
 		default: edge_mask_reg_512p3[135] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b10001010001,
13'b10001010010,
13'b10001010011,
13'b10001010100,
13'b10001010101,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010101000,
13'b10010101001,
13'b11001000000,
13'b11001000001,
13'b11001000010,
13'b11001000011,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001010000,
13'b11001010001,
13'b11001010010,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100010,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b100000110000,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001000000,
13'b100001000001,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010000,
13'b100001010001,
13'b100001010010,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110011,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001111000,
13'b110001111001,
13'b110010001000,
13'b110010001001,
13'b111000010010,
13'b111000010011,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000101000,
13'b111000101001,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000111000,
13'b111000111001,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001001000,
13'b111001001001,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001011000,
13'b111001011001,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b1000000100011,
13'b1000000100100,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001100011,
13'b1000001100100,
13'b1000001110011,
13'b1000001110100,
13'b1001000110011,
13'b1001000110100,
13'b1001001000011,
13'b1001001000100,
13'b1001001010011,
13'b1001001010100,
13'b1001001100011,
13'b1001001100100: edge_mask_reg_512p3[136] <= 1'b1;
 		default: edge_mask_reg_512p3[136] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100111,
13'b11010101000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100111,
13'b100010101000,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100111,
13'b101010101000,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010000,
13'b110001010001,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100000,
13'b110001100001,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110001,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010111,
13'b110010011000,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b1000000100100,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1001000100011,
13'b1001000100100,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1010000100010,
13'b1010000100011,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001110000,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1011000100010,
13'b1011000110010,
13'b1011000110011,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001010000,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001100000,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001110010,
13'b1011001110011,
13'b1100001000010,
13'b1100001000011,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1100001100010,
13'b1100001100011: edge_mask_reg_512p3[137] <= 1'b1;
 		default: edge_mask_reg_512p3[137] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010111,
13'b110010011000,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110100,
13'b111001110101,
13'b1000000100100,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1001000100011,
13'b1001000100100,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1010000100010,
13'b1010000100011,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001110000,
13'b1010001110010,
13'b1010001110011,
13'b1011000100010,
13'b1011000110010,
13'b1011000110011,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001010000,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001100000,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1100001000010,
13'b1100001000011,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1100001100010,
13'b1100001100011: edge_mask_reg_512p3[138] <= 1'b1;
 		default: edge_mask_reg_512p3[138] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b1000000100100,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1001000100011,
13'b1001000100100,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1010000100010,
13'b1010000100011,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001110000,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010010000000,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010010000,
13'b1010010010001,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1011000100010,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001010000,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001100000,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001110000,
13'b1011001110001,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011010000000,
13'b1011010000001,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010010000,
13'b1011010010001,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010100001,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1100001000010,
13'b1100001000011,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1100001100000,
13'b1100001100001,
13'b1100001100010,
13'b1100001100011,
13'b1100001100100,
13'b1100001110000,
13'b1100001110001,
13'b1100001110010,
13'b1100001110011,
13'b1100001110100,
13'b1100010000000,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010000,
13'b1100010010001,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010100001,
13'b1100010100010,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010110001,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1101001100000,
13'b1101001100001,
13'b1101001100010,
13'b1101001100011,
13'b1101001110000,
13'b1101001110001,
13'b1101001110010,
13'b1101001110011,
13'b1101001110100,
13'b1101010000000,
13'b1101010000001,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010010001,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010100001,
13'b1101010100010,
13'b1101010100011,
13'b1101010100100,
13'b1101010110001,
13'b1101010110010,
13'b1101010110011,
13'b1101010110100,
13'b1110010000001,
13'b1110010000011,
13'b1110010000100,
13'b1110010010001,
13'b1110010010010,
13'b1110010010011,
13'b1110010010100,
13'b1110010100001,
13'b1110010100010,
13'b1110010100011,
13'b1110010100100,
13'b1110010110011,
13'b1110010110100: edge_mask_reg_512p3[139] <= 1'b1;
 		default: edge_mask_reg_512p3[139] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000110,
13'b100100000111,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110110,
13'b110011110111,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b1000000100100,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1000011010100,
13'b1001000100011,
13'b1001000100100,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001010000000,
13'b1001010000001,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010010000,
13'b1001010010001,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100000,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110000,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1010000100010,
13'b1010000100011,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001110000,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010010000000,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010010000,
13'b1010010010001,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010100000,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110000,
13'b1010010110001,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000000,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1011000100010,
13'b1011000110010,
13'b1011000110011,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001010000,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001100000,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001110000,
13'b1011001110001,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011010000000,
13'b1011010000001,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010010000,
13'b1011010010001,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010100000,
13'b1011010100001,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010110000,
13'b1011010110001,
13'b1011010110010,
13'b1011010110011,
13'b1011010110100,
13'b1011011000000,
13'b1011011000001,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1011011010010,
13'b1011011010011,
13'b1100001000010,
13'b1100001000011,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1100001100000,
13'b1100001100001,
13'b1100001100010,
13'b1100001100011,
13'b1100001110000,
13'b1100001110001,
13'b1100001110010,
13'b1100001110011,
13'b1100010000000,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010010000,
13'b1100010010001,
13'b1100010010010,
13'b1100010010011,
13'b1100010100000,
13'b1100010100001,
13'b1100010100010,
13'b1100010100011,
13'b1100010110000,
13'b1100010110001,
13'b1100010110010,
13'b1100010110011,
13'b1100011000000,
13'b1100011000001,
13'b1100011000010,
13'b1100011000011,
13'b1100011010010,
13'b1100011010011: edge_mask_reg_512p3[140] <= 1'b1;
 		default: edge_mask_reg_512p3[140] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[141] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[142] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000110,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110110,
13'b110001110111,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010100,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000010111,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010011,
13'b1001001010100,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000000110,
13'b1010000000111,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000010111,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001010011,
13'b1010001010100,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000000101,
13'b1011000000110,
13'b1011000000111,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000010110,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001010011,
13'b1100000000010,
13'b1100000000011,
13'b1100000000100,
13'b1100000000101,
13'b1100000000110,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000010100,
13'b1100000010101,
13'b1100000010110,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1100001000011,
13'b1100001000100,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000000100,
13'b1101000000101,
13'b1101000000110,
13'b1101000010001,
13'b1101000010010,
13'b1101000010011,
13'b1101000010100,
13'b1101000010101,
13'b1101000010110,
13'b1101000100000,
13'b1101000100001,
13'b1101000100010,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000110000,
13'b1101000110001,
13'b1101000110010,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101001000000,
13'b1101001000001,
13'b1101001000010,
13'b1101001000011,
13'b1101001000100,
13'b1101001010000,
13'b1101001010010,
13'b1110000000001,
13'b1110000000010,
13'b1110000000011,
13'b1110000000100,
13'b1110000000101,
13'b1110000000110,
13'b1110000010001,
13'b1110000010010,
13'b1110000010011,
13'b1110000010100,
13'b1110000010101,
13'b1110000010110,
13'b1110000100000,
13'b1110000100001,
13'b1110000100010,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000110000,
13'b1110000110001,
13'b1110000110010,
13'b1110000110011,
13'b1110000110100,
13'b1110001000000,
13'b1110001000001,
13'b1110001000010,
13'b1110001000011,
13'b1110001000100,
13'b1111000000010,
13'b1111000000011,
13'b1111000000100,
13'b1111000000101,
13'b1111000000110,
13'b1111000010001,
13'b1111000010010,
13'b1111000010011,
13'b1111000010100,
13'b1111000010101,
13'b1111000100001,
13'b1111000100010,
13'b1111000100011,
13'b1111000110001,
13'b1111000110010: edge_mask_reg_512p3[143] <= 1'b1;
 		default: edge_mask_reg_512p3[143] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000110,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110110,
13'b110001110111,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010100,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010011,
13'b1001001010100,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000000110,
13'b1010000000111,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001010011,
13'b1010001010100,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000000101,
13'b1011000000110,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000010110,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001010011,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000000100,
13'b1100000000101,
13'b1100000000110,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000010100,
13'b1100000010101,
13'b1100000010110,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1100001000011,
13'b1100001000100,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000000100,
13'b1101000000101,
13'b1101000000110,
13'b1101000010001,
13'b1101000010010,
13'b1101000010011,
13'b1101000010100,
13'b1101000010101,
13'b1101000100000,
13'b1101000100001,
13'b1101000100010,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000110000,
13'b1101000110001,
13'b1101000110010,
13'b1101000110011,
13'b1101000110100,
13'b1101001000000,
13'b1101001000001,
13'b1101001000010,
13'b1101001000011,
13'b1101001000100,
13'b1101001010000,
13'b1101001010010,
13'b1110000000001,
13'b1110000000010,
13'b1110000000011,
13'b1110000000100,
13'b1110000000101,
13'b1110000000110,
13'b1110000010001,
13'b1110000010010,
13'b1110000010011,
13'b1110000010100,
13'b1110000010101,
13'b1110000100000,
13'b1110000100001,
13'b1110000100010,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000110000,
13'b1110000110001,
13'b1110000110010,
13'b1110000110011,
13'b1110000110100,
13'b1110001000000,
13'b1110001000001,
13'b1110001000010,
13'b1110001000011,
13'b1111000000001,
13'b1111000000010,
13'b1111000000011,
13'b1111000000100,
13'b1111000000101,
13'b1111000010001,
13'b1111000010010,
13'b1111000010011,
13'b1111000010100,
13'b1111000010101,
13'b1111000100001,
13'b1111000100010: edge_mask_reg_512p3[144] <= 1'b1;
 		default: edge_mask_reg_512p3[144] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000100,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010100,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100100,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000100,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010100,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100100,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110100,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b10010100101,
13'b10010100110,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11110000100,
13'b11110000101,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100110000100,
13'b100110000101,
13'b101010110101,
13'b101010110110,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101110100,
13'b101101110101,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101100100,
13'b110101100101,
13'b111011100100,
13'b111011100101,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101010010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101010001,
13'b1000101010010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101010001,
13'b1001101010010,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100100000,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101010000,
13'b1011101010001,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011110001,
13'b1100011110010,
13'b1100011110011,
13'b1100011110100,
13'b1100100000000,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100000100,
13'b1100100010000,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100000,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101010000,
13'b1100101010001,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011110001,
13'b1101011110010,
13'b1101011110011,
13'b1101011110100,
13'b1101100000000,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100000100,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100010100,
13'b1101100100000,
13'b1101100100001,
13'b1101100100010,
13'b1101100100011,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1110011100010,
13'b1110011100011,
13'b1110011110000,
13'b1110011110001,
13'b1110011110010,
13'b1110011110011,
13'b1110011110100,
13'b1110100000000,
13'b1110100000001,
13'b1110100000010,
13'b1110100000011,
13'b1110100000100,
13'b1110100010000,
13'b1110100010001,
13'b1110100010010,
13'b1110100010011,
13'b1110100010100,
13'b1110100100000,
13'b1110100100001,
13'b1110100100010,
13'b1110100100011,
13'b1110100110000,
13'b1111011110000,
13'b1111011110001,
13'b1111011110010,
13'b1111011110011,
13'b1111100000000,
13'b1111100000001,
13'b1111100000010,
13'b1111100000011,
13'b1111100010000,
13'b1111100010001,
13'b1111100010010,
13'b1111100100000,
13'b1111100100001,
13'b1111100110000: edge_mask_reg_512p3[145] <= 1'b1;
 		default: edge_mask_reg_512p3[145] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100100,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010100,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010100,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100100,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110100,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b10010100101,
13'b10010100110,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110100100,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110100100,
13'b11110100101,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110100100,
13'b100110100101,
13'b101010110101,
13'b101010110110,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010100,
13'b101110010101,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110100,
13'b110101110101,
13'b110110000100,
13'b110110000101,
13'b111011100100,
13'b111011100101,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100100000,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101100000,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011110001,
13'b1100011110010,
13'b1100011110011,
13'b1100011110100,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100000100,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100000,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101100000,
13'b1100101100001,
13'b1100101100010,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011110001,
13'b1101011110010,
13'b1101011110011,
13'b1101011110100,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100000100,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100010100,
13'b1101100100000,
13'b1101100100001,
13'b1101100100010,
13'b1101100100011,
13'b1101100100100,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1110011100010,
13'b1110011100011,
13'b1110011110001,
13'b1110011110010,
13'b1110011110011,
13'b1110011110100,
13'b1110100000000,
13'b1110100000001,
13'b1110100000010,
13'b1110100000011,
13'b1110100000100,
13'b1110100010000,
13'b1110100010001,
13'b1110100010010,
13'b1110100010011,
13'b1110100010100,
13'b1110100100000,
13'b1110100100001,
13'b1110100100010,
13'b1110100100011,
13'b1110100110000,
13'b1110100110001,
13'b1110100110010,
13'b1110100110011,
13'b1110101000000,
13'b1110101000001,
13'b1110101000010,
13'b1110101010000,
13'b1110101010001,
13'b1110101100000,
13'b1111011110000,
13'b1111011110001,
13'b1111011110010,
13'b1111011110011,
13'b1111100000000,
13'b1111100000001,
13'b1111100000010,
13'b1111100000011,
13'b1111100010000,
13'b1111100010001,
13'b1111100010010,
13'b1111100100000,
13'b1111100100001,
13'b1111100100010,
13'b1111100110000,
13'b1111100110001,
13'b1111100110010,
13'b1111101000000,
13'b1111101000001,
13'b1111101010000,
13'b1111101010001: edge_mask_reg_512p3[146] <= 1'b1;
 		default: edge_mask_reg_512p3[146] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b10010100101,
13'b10010100110,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010101,
13'b11101010110,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101010101,
13'b100101010110,
13'b101010110101,
13'b101010110110,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101010101,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000101,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100010,
13'b1000100100011,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100010,
13'b1001100100011,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100010,
13'b1010100100011,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1100011100001,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011110000,
13'b1100011110001,
13'b1100011110010,
13'b1100011110011,
13'b1100011110100,
13'b1100100000000,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100000100,
13'b1100100010000,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100001,
13'b1100100100010,
13'b1101011100001,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011110000,
13'b1101011110001,
13'b1101011110010,
13'b1101011110011,
13'b1101011110100,
13'b1101100000000,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100000100,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100010100,
13'b1101100100001,
13'b1101100100010,
13'b1110011100010,
13'b1110011100011,
13'b1110011110000,
13'b1110011110001,
13'b1110011110010,
13'b1110011110011,
13'b1110011110100,
13'b1110100000000,
13'b1110100000001,
13'b1110100000010,
13'b1110100000011,
13'b1110100000100,
13'b1110100010000,
13'b1110100010001,
13'b1110100010010,
13'b1110100010011,
13'b1110100010100,
13'b1111011110000,
13'b1111011110001,
13'b1111011110010,
13'b1111011110011,
13'b1111100000000,
13'b1111100000001,
13'b1111100000010,
13'b1111100000011,
13'b1111100010000,
13'b1111100010001,
13'b1111100010010: edge_mask_reg_512p3[147] <= 1'b1;
 		default: edge_mask_reg_512p3[147] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b100001110110,
13'b100001110111,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b101001110110,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b111010100101,
13'b111010100110,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100010100,
13'b111100010101,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011011110101,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100010011,
13'b1011100010100,
13'b1100010100100,
13'b1100010100101,
13'b1100010110011,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100011000011,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011010010,
13'b1100011010011,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011100101,
13'b1100011110010,
13'b1100011110011,
13'b1100011110100,
13'b1100011110101,
13'b1100100000010,
13'b1100100000011,
13'b1100100000100,
13'b1100100000101,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1101010100100,
13'b1101010100101,
13'b1101010110011,
13'b1101010110100,
13'b1101010110101,
13'b1101011000011,
13'b1101011000100,
13'b1101011000101,
13'b1101011010010,
13'b1101011010011,
13'b1101011010100,
13'b1101011010101,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011100101,
13'b1101011110010,
13'b1101011110011,
13'b1101011110100,
13'b1101011110101,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100000100,
13'b1101100010010,
13'b1101100010011,
13'b1101100010100,
13'b1110010100100,
13'b1110010100101,
13'b1110010110011,
13'b1110010110100,
13'b1110010110101,
13'b1110011000010,
13'b1110011000011,
13'b1110011000100,
13'b1110011000101,
13'b1110011010010,
13'b1110011010011,
13'b1110011010100,
13'b1110011010101,
13'b1110011100001,
13'b1110011100010,
13'b1110011100011,
13'b1110011100100,
13'b1110011100101,
13'b1110011110001,
13'b1110011110010,
13'b1110011110011,
13'b1110011110100,
13'b1110011110101,
13'b1110100000001,
13'b1110100000010,
13'b1110100000011,
13'b1110100000100,
13'b1110100010010,
13'b1110100010011,
13'b1110100010100,
13'b1111010100100,
13'b1111010100101,
13'b1111010110010,
13'b1111010110011,
13'b1111010110100,
13'b1111010110101,
13'b1111011000001,
13'b1111011000010,
13'b1111011000011,
13'b1111011000100,
13'b1111011000101,
13'b1111011010001,
13'b1111011010010,
13'b1111011010011,
13'b1111011010100,
13'b1111011010101,
13'b1111011100001,
13'b1111011100010,
13'b1111011100011,
13'b1111011100100,
13'b1111011100101,
13'b1111011110001,
13'b1111011110010,
13'b1111011110011,
13'b1111011110100,
13'b1111100000001,
13'b1111100000010,
13'b1111100000011: edge_mask_reg_512p3[148] <= 1'b1;
 		default: edge_mask_reg_512p3[148] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b100001100101,
13'b100001100110,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b101001100101,
13'b101001100110,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b110001110101,
13'b110001110110,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b111010010100,
13'b111010010101,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100010100,
13'b111100010101,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1010010010011,
13'b1010010010100,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010110010,
13'b1011010110011,
13'b1011010110100,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1011011010010,
13'b1011011010011,
13'b1011011010100,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010011,
13'b1011100010100,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010100010,
13'b1100010100011,
13'b1100010100100,
13'b1100010110001,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100011000001,
13'b1100011000010,
13'b1100011000011,
13'b1100011000100,
13'b1100011010010,
13'b1100011010011,
13'b1100011010100,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011110010,
13'b1100011110011,
13'b1100011110100,
13'b1100100000010,
13'b1100100000011,
13'b1100100000100,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1101010010010,
13'b1101010010011,
13'b1101010100001,
13'b1101010100010,
13'b1101010100011,
13'b1101010100100,
13'b1101010110001,
13'b1101010110010,
13'b1101010110011,
13'b1101010110100,
13'b1101011000001,
13'b1101011000010,
13'b1101011000011,
13'b1101011000100,
13'b1101011010001,
13'b1101011010010,
13'b1101011010011,
13'b1101011010100,
13'b1101011100001,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011110001,
13'b1101011110010,
13'b1101011110011,
13'b1101011110100,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100000100,
13'b1101100010010,
13'b1101100010011,
13'b1101100010100,
13'b1110010010010,
13'b1110010010011,
13'b1110010100000,
13'b1110010100001,
13'b1110010100010,
13'b1110010100011,
13'b1110010110000,
13'b1110010110001,
13'b1110010110010,
13'b1110010110011,
13'b1110010110100,
13'b1110011000000,
13'b1110011000001,
13'b1110011000010,
13'b1110011000011,
13'b1110011000100,
13'b1110011010000,
13'b1110011010001,
13'b1110011010010,
13'b1110011010011,
13'b1110011010100,
13'b1110011100000,
13'b1110011100001,
13'b1110011100010,
13'b1110011100011,
13'b1110011100100,
13'b1110011110000,
13'b1110011110001,
13'b1110011110010,
13'b1110011110011,
13'b1110011110100,
13'b1110100000001,
13'b1110100000010,
13'b1110100000011,
13'b1110100000100,
13'b1110100010010,
13'b1110100010011,
13'b1110100010100,
13'b1111010100000,
13'b1111010100001,
13'b1111010100010,
13'b1111010110000,
13'b1111010110001,
13'b1111010110010,
13'b1111011000000,
13'b1111011000001,
13'b1111011000010,
13'b1111011000011,
13'b1111011010000,
13'b1111011010001,
13'b1111011010010,
13'b1111011010011,
13'b1111011100000,
13'b1111011100001,
13'b1111011100010,
13'b1111011100011,
13'b1111011110000,
13'b1111011110001,
13'b1111011110010,
13'b1111011110011,
13'b1111100000000,
13'b1111100000001,
13'b1111100000010,
13'b1111100000011: edge_mask_reg_512p3[149] <= 1'b1;
 		default: edge_mask_reg_512p3[149] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10010100101,
13'b10010100110,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b101010110101,
13'b101010110110,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b111011100100,
13'b111011100101,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100011,
13'b1000101100100,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011110010,
13'b1100011110011,
13'b1100011110100,
13'b1100100000010,
13'b1100100000011,
13'b1100100000100,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011110001,
13'b1101011110010,
13'b1101011110011,
13'b1101011110100,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100000100,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100010100,
13'b1101100100000,
13'b1101100100001,
13'b1101100100010,
13'b1101100100011,
13'b1101100100100,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101100110100,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1110011100010,
13'b1110011100011,
13'b1110011110001,
13'b1110011110010,
13'b1110011110011,
13'b1110011110100,
13'b1110100000000,
13'b1110100000001,
13'b1110100000010,
13'b1110100000011,
13'b1110100000100,
13'b1110100010000,
13'b1110100010001,
13'b1110100010010,
13'b1110100010011,
13'b1110100010100,
13'b1110100100000,
13'b1110100100001,
13'b1110100100010,
13'b1110100100011,
13'b1110100100100,
13'b1110100110000,
13'b1110100110001,
13'b1110100110010,
13'b1110100110011,
13'b1110101000000,
13'b1110101000001,
13'b1110101000010,
13'b1110101000011,
13'b1110101010000,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101100000,
13'b1110101100010,
13'b1111011110000,
13'b1111011110001,
13'b1111011110010,
13'b1111011110011,
13'b1111100000000,
13'b1111100000001,
13'b1111100000010,
13'b1111100000011,
13'b1111100010000,
13'b1111100010001,
13'b1111100010010,
13'b1111100010011,
13'b1111100100000,
13'b1111100100001,
13'b1111100100010,
13'b1111100110000,
13'b1111100110001,
13'b1111100110010,
13'b1111101000000,
13'b1111101000001,
13'b1111101000010,
13'b1111101010000,
13'b1111101010001: edge_mask_reg_512p3[150] <= 1'b1;
 		default: edge_mask_reg_512p3[150] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[151] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100111,
13'b1001101000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b111000010111,
13'b111000011000,
13'b111000100111,
13'b111000101000,
13'b1000000010111,
13'b1000000011000,
13'b1000000100111,
13'b1000000101000,
13'b1001000010110,
13'b1001000010111,
13'b1001000011000,
13'b1001000100111,
13'b1001000101000,
13'b1010000000110,
13'b1010000000111,
13'b1010000001000,
13'b1010000010110,
13'b1010000010111,
13'b1010000011000,
13'b1010000100111,
13'b1010000101000,
13'b1011000000110,
13'b1011000000111,
13'b1011000001000,
13'b1011000010110,
13'b1011000010111,
13'b1011000011000,
13'b1011000100111,
13'b1011000101000,
13'b1100000000110,
13'b1100000000111,
13'b1100000001000,
13'b1100000010110,
13'b1100000010111,
13'b1100000011000,
13'b1100000100111,
13'b1100000101000,
13'b1101000000110,
13'b1101000000111,
13'b1101000001000,
13'b1101000010110,
13'b1101000010111,
13'b1101000011000,
13'b1101000100110,
13'b1101000100111,
13'b1101000101000,
13'b1110000000110,
13'b1110000000111,
13'b1110000001000,
13'b1110000010110,
13'b1110000010111,
13'b1110000011000,
13'b1110000100110,
13'b1110000100111,
13'b1110000101000,
13'b1111000000110,
13'b1111000000111,
13'b1111000001000,
13'b1111000010110,
13'b1111000010111,
13'b1111000011000,
13'b1111000100111,
13'b1111000101000: edge_mask_reg_512p3[152] <= 1'b1;
 		default: edge_mask_reg_512p3[152] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[153] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000110,
13'b100001000111,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000110,
13'b101001000111,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110110,
13'b110000110111,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010010,
13'b1100000010011,
13'b1101000000000,
13'b1101000000001: edge_mask_reg_512p3[154] <= 1'b1;
 		default: edge_mask_reg_512p3[154] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000101,
13'b11001000110,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100001000101,
13'b100001000110,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110101,
13'b101000110110,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000110101,
13'b111000010000: edge_mask_reg_512p3[155] <= 1'b1;
 		default: edge_mask_reg_512p3[155] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000110,
13'b10010000111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000110,
13'b11010000111,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000110,
13'b100010000111,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110110,
13'b110001110111,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1101000000000,
13'b1101000000001,
13'b1101000010000,
13'b1101000010001,
13'b1101000100000,
13'b1101000100001,
13'b1101000110000,
13'b1101000110001,
13'b1101001000000,
13'b1101001000001,
13'b1110000000000,
13'b1110000000001,
13'b1110000010000,
13'b1110000010001,
13'b1110000100000,
13'b1110000100001,
13'b1110000110000,
13'b1110000110001,
13'b1110001000000,
13'b1110001000001,
13'b1111000000000,
13'b1111000000001,
13'b1111000010000,
13'b1111000010001,
13'b1111000100000,
13'b1111000100001: edge_mask_reg_512p3[156] <= 1'b1;
 		default: edge_mask_reg_512p3[156] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100000,
13'b11101100001,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110000,
13'b11101110001,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000000,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010000,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100000,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110000,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110100010111,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000111,
13'b111101001000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010111,
13'b111101011000,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100111,
13'b111101101000,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110110,
13'b111110110111,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000110,
13'b111111000111,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b1000101000001,
13'b1000101000010,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111010000,
13'b1000111010001,
13'b1001101100010,
13'b1001101110001,
13'b1001101110010: edge_mask_reg_512p3[157] <= 1'b1;
 		default: edge_mask_reg_512p3[157] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000100101,
13'b101000100110: edge_mask_reg_512p3[158] <= 1'b1;
 		default: edge_mask_reg_512p3[158] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000100101,
13'b101000100110: edge_mask_reg_512p3[159] <= 1'b1;
 		default: edge_mask_reg_512p3[159] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101110011000,
13'b101110011001,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110101000,
13'b110110101001,
13'b110110110110,
13'b110110111000,
13'b110110111001,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110110101,
13'b111110110110,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001110110100,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1011111000100,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111110010,
13'b1100111110011,
13'b1101111010010,
13'b1101111010011,
13'b1101111100010,
13'b1101111100011,
13'b1101111110010,
13'b1101111110011: edge_mask_reg_512p3[160] <= 1'b1;
 		default: edge_mask_reg_512p3[160] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101100111,
13'b100101101000,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101101000,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000010,
13'b110110000011,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110101000,
13'b111110101001,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110111000,
13'b111110111001,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100000,
13'b111111100001,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010110110011,
13'b1010110110100,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111110010,
13'b1100111110011,
13'b1101111010010,
13'b1101111010011,
13'b1101111100010,
13'b1101111100011: edge_mask_reg_512p3[161] <= 1'b1;
 		default: edge_mask_reg_512p3[161] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[162] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[163] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011011000,
13'b110011011001,
13'b111001000111,
13'b111001001000,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011001000,
13'b111011001001,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000001111001,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010001001,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010011010,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010101010,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1001001000110,
13'b1001001000111,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001001111001,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010001001,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010011010,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010101010,
13'b1001010111000,
13'b1001010111001,
13'b1001010111010,
13'b1001011001000,
13'b1001011001001,
13'b1010001000111,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1010001100110,
13'b1010001100111,
13'b1010001101000,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010001111001,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010001001,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010011010,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010101010,
13'b1010010111000,
13'b1010010111001,
13'b1010010111010,
13'b1010011001000,
13'b1010011001001,
13'b1011001000110,
13'b1011001000111,
13'b1011001010101,
13'b1011001010110,
13'b1011001010111,
13'b1011001011000,
13'b1011001100110,
13'b1011001100111,
13'b1011001101000,
13'b1011001110110,
13'b1011001110111,
13'b1011001111000,
13'b1011001111001,
13'b1011010000110,
13'b1011010000111,
13'b1011010001000,
13'b1011010001001,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010011001,
13'b1011010011010,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010101010,
13'b1011010111000,
13'b1011010111001,
13'b1011010111010,
13'b1011011001000,
13'b1011011001001,
13'b1100001000101,
13'b1100001000110,
13'b1100001010101,
13'b1100001010110,
13'b1100001010111,
13'b1100001100101,
13'b1100001100110,
13'b1100001100111,
13'b1100001101000,
13'b1100001110101,
13'b1100001110110,
13'b1100001110111,
13'b1100001111000,
13'b1100001111001,
13'b1100010000110,
13'b1100010000111,
13'b1100010001000,
13'b1100010001001,
13'b1100010010110,
13'b1100010010111,
13'b1100010011000,
13'b1100010011001,
13'b1100010011010,
13'b1100010100111,
13'b1100010101000,
13'b1100010101001,
13'b1100010101010,
13'b1100010111000,
13'b1100010111001,
13'b1100010111010,
13'b1100011001001,
13'b1100011001010,
13'b1101001000110,
13'b1101001010100,
13'b1101001010101,
13'b1101001010110,
13'b1101001010111,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001100110,
13'b1101001100111,
13'b1101001101000,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101001110110,
13'b1101001110111,
13'b1101001111000,
13'b1101001111001,
13'b1101010000101,
13'b1101010000110,
13'b1101010000111,
13'b1101010001000,
13'b1101010001001,
13'b1101010001010,
13'b1101010010110,
13'b1101010010111,
13'b1101010011000,
13'b1101010011001,
13'b1101010011010,
13'b1101010100111,
13'b1101010101000,
13'b1101010101001,
13'b1101010101010,
13'b1101010111000,
13'b1101010111001,
13'b1101010111010,
13'b1101011001001,
13'b1101011001010,
13'b1110001000110,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001010110,
13'b1110001010111,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001100110,
13'b1110001100111,
13'b1110001101000,
13'b1110001110011,
13'b1110001110100,
13'b1110001110101,
13'b1110001110110,
13'b1110001110111,
13'b1110001111000,
13'b1110001111001,
13'b1110010000100,
13'b1110010000101,
13'b1110010000110,
13'b1110010000111,
13'b1110010001000,
13'b1110010001001,
13'b1110010001010,
13'b1110010010101,
13'b1110010010110,
13'b1110010010111,
13'b1110010011000,
13'b1110010011001,
13'b1110010011010,
13'b1110010100110,
13'b1110010100111,
13'b1110010101000,
13'b1110010101001,
13'b1110010101010,
13'b1110010110111,
13'b1110010111000,
13'b1110010111001,
13'b1110010111010,
13'b1110011001001,
13'b1111001010101,
13'b1111001010110,
13'b1111001010111,
13'b1111001100011,
13'b1111001100100,
13'b1111001100101,
13'b1111001100110,
13'b1111001100111,
13'b1111001101000,
13'b1111001110011,
13'b1111001110100,
13'b1111001110101,
13'b1111001110110,
13'b1111001110111,
13'b1111001111000,
13'b1111010000100,
13'b1111010000101,
13'b1111010000110,
13'b1111010000111,
13'b1111010001000,
13'b1111010001001,
13'b1111010010101,
13'b1111010010110,
13'b1111010010111,
13'b1111010011000,
13'b1111010011001,
13'b1111010011010,
13'b1111010100110,
13'b1111010100111,
13'b1111010101000,
13'b1111010101001,
13'b1111010101010,
13'b1111010110111,
13'b1111010111000,
13'b1111010111001,
13'b1111010111010: edge_mask_reg_512p3[164] <= 1'b1;
 		default: edge_mask_reg_512p3[164] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b100000111000,
13'b100000111001,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010110101,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010000,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100000,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000000,
13'b1001010000001,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010000,
13'b1001010010001,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100000,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010010000000,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010010000,
13'b1010010010001,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001110001,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011010000001,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010010001,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010100001,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1100001110100,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010010,
13'b1100010010100,
13'b1100010010101,
13'b1100010100100: edge_mask_reg_512p3[165] <= 1'b1;
 		default: edge_mask_reg_512p3[165] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010111,
13'b100011000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100001000,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100001000,
13'b100000111000,
13'b100000111001,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100001000,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b110001011000,
13'b110001011001,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b111001100101,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010100,
13'b111011010101,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010100,
13'b1000011010101,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000001,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010001,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010010001,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110001,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011010011,
13'b1010011010100,
13'b1011001100100,
13'b1011001100101,
13'b1011001110001,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011010000001,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010010001,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010100001,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010110001,
13'b1011010110010,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011011000001,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1011011010011,
13'b1100001110100,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010001,
13'b1100010010010,
13'b1100010010100,
13'b1100010010101,
13'b1100010100011,
13'b1100010100100,
13'b1100010110011,
13'b1100010110100: edge_mask_reg_512p3[166] <= 1'b1;
 		default: edge_mask_reg_512p3[166] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[167] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000001,
13'b1110000010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010001,
13'b1110010010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100001,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110001,
13'b10101110010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000001,
13'b10110000010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010000,
13'b10110010001,
13'b10110010010,
13'b10110010011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100000,
13'b10110100001,
13'b10110100010,
13'b10110100011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010000,
13'b11101010001,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000000,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110000,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100101000,
13'b100100101001,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100101000,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110111000,
13'b110110111001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111001000,
13'b110111001001,
13'b110111010011,
13'b110111011000,
13'b110111011001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101101000,
13'b111101110010,
13'b111101110011,
13'b111101111000,
13'b111101111001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110001000,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110011000,
13'b111110100010,
13'b111110100011,
13'b111110101000,
13'b111110111000: edge_mask_reg_512p3[168] <= 1'b1;
 		default: edge_mask_reg_512p3[168] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[169] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000110,
13'b10010000111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000110,
13'b11010000111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000110,
13'b100010000111,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110110,
13'b110001110111,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1101000000000,
13'b1101000000001,
13'b1101000010000,
13'b1101000010001,
13'b1101000100000,
13'b1101000100001,
13'b1101000110000,
13'b1101000110001,
13'b1101001000000,
13'b1101001000001,
13'b1110000000000,
13'b1110000000001,
13'b1110000010000,
13'b1110000010001,
13'b1110000100000,
13'b1110000100001,
13'b1110000110000,
13'b1110000110001,
13'b1110001000000,
13'b1110001000001: edge_mask_reg_512p3[170] <= 1'b1;
 		default: edge_mask_reg_512p3[170] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010110,
13'b101010010111,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110011,
13'b110001110100,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000110,
13'b110010000111,
13'b110010010110,
13'b110010010111,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010111,
13'b111000011000,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010111,
13'b111001011000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100111,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001110001,
13'b1001001110010,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001110001: edge_mask_reg_512p3[171] <= 1'b1;
 		default: edge_mask_reg_512p3[171] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110000,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000000,
13'b10010000001,
13'b10010000010,
13'b10010000011,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010000,
13'b10010010001,
13'b10010010010,
13'b10010010011,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100000,
13'b10010100001,
13'b10010100010,
13'b10010100011,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110000,
13'b10010110001,
13'b10010110010,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010000,
13'b11001010001,
13'b11001010010,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100000,
13'b11001100001,
13'b11001100010,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110000,
13'b11001110001,
13'b11001110010,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000000,
13'b11010000001,
13'b11010000010,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010000,
13'b11010010001,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100000,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110000,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000000,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010000,
13'b100001010001,
13'b100001010010,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100000,
13'b100001100001,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110000,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000000,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010000,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100000,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010110000,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100011000000,
13'b100011000001,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101011000000,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011010101,
13'b101011010110,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110000,
13'b110010110001,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000101,
13'b110011000110,
13'b110011010101,
13'b110011010110,
13'b111000100010,
13'b111000100011,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010101,
13'b111010010110,
13'b111010100000,
13'b111010100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010010000,
13'b1000010010001,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001010000000,
13'b1001010000001,
13'b1001010000010,
13'b1010000110001,
13'b1010000110010,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001110001,
13'b1010001110010: edge_mask_reg_512p3[172] <= 1'b1;
 		default: edge_mask_reg_512p3[172] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101001000,
13'b101101001001,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100100,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101100011,
13'b111101100100,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110001000,
13'b111110001001,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110011000,
13'b111110011001,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010111,
13'b111111011000,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100111,
13'b111111101000,
13'b1000101100011,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111100000,
13'b1001111100001,
13'b1010101110001,
13'b1010101110010,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111010000,
13'b1010111010001,
13'b1010111100000,
13'b1011101110001,
13'b1011101110010,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011111000000,
13'b1011111000001,
13'b1100101110010,
13'b1100110000001,
13'b1100110000010,
13'b1100110010001,
13'b1100110010010,
13'b1100110100001,
13'b1100110100010: edge_mask_reg_512p3[173] <= 1'b1;
 		default: edge_mask_reg_512p3[173] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011010,
13'b10011011,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11111000,
13'b11111001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011101001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011101001,
13'b11011101010,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b101000101000,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010111000,
13'b110010111001,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110101,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110101,
13'b1010001010011,
13'b1010001010100,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001110001,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011010000001,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010100101,
13'b1100001100001,
13'b1100001100010,
13'b1100001100011,
13'b1100001110001,
13'b1100001110010,
13'b1100001110011,
13'b1100001110100,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1101001100010,
13'b1101001110010,
13'b1101001110011,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100: edge_mask_reg_512p3[174] <= 1'b1;
 		default: edge_mask_reg_512p3[174] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100101,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010100,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100100,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110100,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b100100000100,
13'b100100000101,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100111000101,
13'b100111000110,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b110100100100,
13'b110100100101,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b111100110011,
13'b111100110100,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b1000100110010,
13'b1000100110011,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1001100110010,
13'b1001100110011,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010011,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110010011,
13'b1011100110001,
13'b1011100110010,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1100100110001,
13'b1100100110010,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1100101110001,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1101100110001,
13'b1101100110010,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1101101110001,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1101110000010,
13'b1101110000011,
13'b1101110000100,
13'b1110101000000,
13'b1110101000001,
13'b1110101000010,
13'b1110101010000,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101100000,
13'b1110101100001,
13'b1110101100010,
13'b1110101100011,
13'b1110101110001,
13'b1110101110010,
13'b1110101110011,
13'b1110110000010,
13'b1110110000011,
13'b1110110000100,
13'b1111101000000,
13'b1111101000001,
13'b1111101010000,
13'b1111101010001,
13'b1111101010010,
13'b1111101100000,
13'b1111101100001,
13'b1111101100010,
13'b1111101100011,
13'b1111101110000,
13'b1111101110001,
13'b1111101110010,
13'b1111101110011,
13'b1111110000010: edge_mask_reg_512p3[175] <= 1'b1;
 		default: edge_mask_reg_512p3[175] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011011,
13'b11011100,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11101101,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b11111101,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100001101,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100011101,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100101101,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b100111101,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101001101,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101011101,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b101101101,
13'b1011101011,
13'b1011101100,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1011111101,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100001101,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100011101,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100101101,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1100111101,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101001101,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101011101,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101101101,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1101111101,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110001101,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b1110011101,
13'b10100001011,
13'b10100001100,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101011101,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101101101,
13'b10101110100,
13'b10101110101,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10101111101,
13'b10110000100,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110001101,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110010100,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111000,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110111,
13'b100110111000,
13'b101100100110,
13'b101100100111,
13'b101100110110,
13'b101100110111,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b110101000110,
13'b110101000111,
13'b110101010110,
13'b110101010111,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110110,
13'b110110110111,
13'b111101010110,
13'b111101010111,
13'b111101100110,
13'b111101100111,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110110,
13'b1000101110110,
13'b1000101110111,
13'b1000110000110,
13'b1000110000111,
13'b1000110010110,
13'b1000110010111,
13'b1000110100110,
13'b1000110100111: edge_mask_reg_512p3[176] <= 1'b1;
 		default: edge_mask_reg_512p3[176] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011100110,
13'b1011100111,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100011110110,
13'b100011110111,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110100000110,
13'b110100000111,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010101,
13'b110111010110,
13'b111100100110,
13'b111100100111,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100101,
13'b111110100110,
13'b111110110101,
13'b111110110110,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100101,
13'b1000110100110,
13'b1000110110101,
13'b1000110110110,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110101,
13'b1001110110110,
13'b1010100100110,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1011100100101,
13'b1011100100110,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1100100100101,
13'b1100100100110,
13'b1100100110101,
13'b1100100110110,
13'b1100101000101,
13'b1100101000110,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100100,
13'b1100101100101,
13'b1100101100110,
13'b1100101110100,
13'b1100101110101,
13'b1100101110110,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110010100,
13'b1100110010101,
13'b1100110010110,
13'b1100110100100,
13'b1100110100101,
13'b1100110100110,
13'b1100110110100,
13'b1100110110101,
13'b1100110110110,
13'b1101100100101,
13'b1101100100110,
13'b1101100110100,
13'b1101100110101,
13'b1101100110110,
13'b1101101000100,
13'b1101101000101,
13'b1101101000110,
13'b1101101010100,
13'b1101101010101,
13'b1101101010110,
13'b1101101100100,
13'b1101101100101,
13'b1101101100110,
13'b1101101110100,
13'b1101101110101,
13'b1101101110110,
13'b1101110000100,
13'b1101110000101,
13'b1101110000110,
13'b1101110010100,
13'b1101110010101,
13'b1101110010110,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1101110110100,
13'b1101110110101,
13'b1101110110110,
13'b1110100100101,
13'b1110100100110,
13'b1110100110100,
13'b1110100110101,
13'b1110100110110,
13'b1110101000100,
13'b1110101000101,
13'b1110101000110,
13'b1110101010100,
13'b1110101010101,
13'b1110101010110,
13'b1110101100100,
13'b1110101100101,
13'b1110101100110,
13'b1110101110100,
13'b1110101110101,
13'b1110101110110,
13'b1110110000100,
13'b1110110000101,
13'b1110110000110,
13'b1110110010100,
13'b1110110010101,
13'b1110110010110,
13'b1110110100100,
13'b1110110100101,
13'b1110110100110,
13'b1110110110100,
13'b1110110110101,
13'b1110110110110,
13'b1111100110101,
13'b1111100110110,
13'b1111101000100,
13'b1111101000101,
13'b1111101000110,
13'b1111101010100,
13'b1111101010101,
13'b1111101010110,
13'b1111101100100,
13'b1111101100101,
13'b1111101100110,
13'b1111101110100,
13'b1111101110101,
13'b1111101110110,
13'b1111110000100,
13'b1111110000101,
13'b1111110000110,
13'b1111110010100,
13'b1111110010101,
13'b1111110010110,
13'b1111110100100,
13'b1111110100101,
13'b1111110100110,
13'b1111110110101,
13'b1111110110110: edge_mask_reg_512p3[177] <= 1'b1;
 		default: edge_mask_reg_512p3[177] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100000,
13'b10100001,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110000,
13'b10110001,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000000,
13'b11000001,
13'b11000010,
13'b11000011,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010000,
13'b11010001,
13'b11010010,
13'b11010011,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100000,
13'b11100001,
13'b11100010,
13'b11100011,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110000,
13'b11110001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010010,
13'b1010010011,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100000,
13'b1010100001,
13'b1010100010,
13'b1010100011,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110000,
13'b1010110001,
13'b1010110010,
13'b1010110011,
13'b1010110100,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000000,
13'b1011000001,
13'b1011000010,
13'b1011000011,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010000,
13'b1011010001,
13'b1011010010,
13'b1011010011,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100000,
13'b1011100001,
13'b1011100010,
13'b1011100011,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110000,
13'b1011110001,
13'b1011110010,
13'b1011110011,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000000,
13'b1100000001,
13'b1100000010,
13'b1100000011,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010000,
13'b1100010001,
13'b1100010010,
13'b1100010011,
13'b1100010100,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100000,
13'b1100100010,
13'b1100100011,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b10001110111,
13'b10001111000,
13'b10010000010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010010,
13'b10010010011,
13'b10010010100,
13'b10010010101,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100000,
13'b10010100001,
13'b10010100010,
13'b10010100011,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110000,
13'b10010110001,
13'b10010110010,
13'b10010110011,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000000,
13'b10011000001,
13'b10011000010,
13'b10011000011,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010000,
13'b10011010001,
13'b10011010010,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100000,
13'b10011100001,
13'b10011100010,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110000,
13'b10011110001,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000000,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010000,
13'b10100010001,
13'b10100010010,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100000,
13'b10100100001,
13'b10100100010,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110000,
13'b10100110001,
13'b10100110010,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000010,
13'b10101000011,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110000,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000000,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010000,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100000,
13'b11011100001,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110000,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000000,
13'b11100000001,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010000,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100000,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110000,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101101000,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110000,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000000,
13'b100100000001,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010000,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100000,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100111,
13'b100101101000,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010111,
13'b101101011000,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101011000,
13'b111011000111,
13'b111011001000,
13'b111011010111,
13'b111011011000,
13'b111011100111,
13'b111011101000,
13'b111011110111,
13'b111011111000,
13'b111100000111,
13'b111100001000,
13'b111100010111,
13'b111100011000,
13'b111100101000: edge_mask_reg_512p3[178] <= 1'b1;
 		default: edge_mask_reg_512p3[178] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011011,
13'b10011100,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11011101,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11101101,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b11111101,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100001101,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100011101,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100101101,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b100111101,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101001101,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101011101,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b101101101,
13'b1010101011,
13'b1010101100,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011101101,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1011111101,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100001101,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100011101,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100101101,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1100111101,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101001101,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101011101,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101101101,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1101111101,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110001101,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b1110011101,
13'b10010111011,
13'b10010111100,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100101101,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10100111101,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101001101,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101011101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101101101,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101011,
13'b10110101100,
13'b11011011011,
13'b11011011100,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111011,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001011,
13'b11100001100,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b111100010100,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000111,
13'b111110001000,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1001101000101,
13'b1001101000110,
13'b1001101010101,
13'b1001101010110,
13'b1001101100101,
13'b1001101100110,
13'b1001101110101,
13'b1001101110110: edge_mask_reg_512p3[179] <= 1'b1;
 		default: edge_mask_reg_512p3[179] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110111,
13'b100111000,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010000,
13'b11011010001,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100000,
13'b11011100001,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110000,
13'b11011110001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000001,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010001,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100101000,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110000,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000000,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010000,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100000,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110000,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000000,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110000,
13'b100011110001,
13'b100011110010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000000,
13'b100100000001,
13'b100100000010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100101000,
13'b100100101001,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000000,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110000,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000000,
13'b101100000001,
13'b101100000010,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010000,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000001,
13'b110100000010,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001101000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001111000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010001000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010011000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101000,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010111000,
13'b111010111001,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011001000,
13'b111011001001,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011011000,
13'b111011011001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011101000,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b1000001010010,
13'b1000001010011,
13'b1000001100010,
13'b1000001100011,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100010,
13'b1000011100011,
13'b1000011110010,
13'b1001001100011,
13'b1001001110010,
13'b1001001110011,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010010010,
13'b1001010010011,
13'b1001010100010,
13'b1001010100011,
13'b1001010110010,
13'b1001010110011,
13'b1001011000010,
13'b1001011000011: edge_mask_reg_512p3[180] <= 1'b1;
 		default: edge_mask_reg_512p3[180] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000111,
13'b101001000,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101101000,
13'b100101101001,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110011,
13'b1010111110100,
13'b1011110010100,
13'b1011110010101,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111110011,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1101110100011,
13'b1101110100100,
13'b1101110100101,
13'b1101110110011,
13'b1101110110100,
13'b1101110110101,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111010011,
13'b1101111010100,
13'b1110110100011,
13'b1110110100100,
13'b1110110100101,
13'b1110110110011,
13'b1110110110100,
13'b1110110110101,
13'b1110111000010,
13'b1110111000011,
13'b1110111000100,
13'b1110111000101,
13'b1110111010011,
13'b1110111010100,
13'b1111110100011,
13'b1111110100100,
13'b1111110100101,
13'b1111110110011,
13'b1111110110100,
13'b1111110110101,
13'b1111111000011,
13'b1111111000100,
13'b1111111000101,
13'b1111111010011,
13'b1111111010100: edge_mask_reg_512p3[181] <= 1'b1;
 		default: edge_mask_reg_512p3[181] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101101001000,
13'b101101001001,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101011000,
13'b110101011001,
13'b110101101000,
13'b110101101001,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111001000,
13'b110111001001,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110011001,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110011001,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110101001,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110010,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010110111000,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011101110111,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110110010,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1100101110101,
13'b1100101110110,
13'b1100101110111,
13'b1100110000001,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110000111,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110100110,
13'b1100110100111,
13'b1100110101000,
13'b1100110110010,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1101110000010,
13'b1101110000011,
13'b1101110000100,
13'b1101110000101,
13'b1101110000110,
13'b1101110000111,
13'b1101110010010,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1101110010110,
13'b1101110010111,
13'b1101110100010,
13'b1101110100011,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1101110100111,
13'b1101110101000,
13'b1101110110110,
13'b1101110110111,
13'b1110110000011,
13'b1110110000100,
13'b1110110000101,
13'b1110110000110,
13'b1110110010011,
13'b1110110010100,
13'b1110110010101,
13'b1110110010110,
13'b1110110100011,
13'b1110110100100,
13'b1110110100101,
13'b1110110100110,
13'b1111110000100,
13'b1111110000101,
13'b1111110010100,
13'b1111110010101,
13'b1111110010110,
13'b1111110100100,
13'b1111110100101,
13'b1111110100110: edge_mask_reg_512p3[182] <= 1'b1;
 		default: edge_mask_reg_512p3[182] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110110,
13'b11011110111,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110110,
13'b100011110111,
13'b101001000110,
13'b101001000111,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110110,
13'b101011110111,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100110,
13'b110011100111,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000100,
13'b1010011000101,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010000110,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010010110,
13'b1100010100001,
13'b1100010100010,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010110001,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100011000011,
13'b1100011000100,
13'b1101001110100,
13'b1101001110101,
13'b1101001110110,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1101010000110,
13'b1101010010001,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010010101,
13'b1101010010110,
13'b1101010100001,
13'b1101010100010,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010100110,
13'b1101010110001,
13'b1101010110010,
13'b1101010110011,
13'b1101010110100,
13'b1101010110101,
13'b1101011000011,
13'b1101011000100,
13'b1110001110100,
13'b1110001110101,
13'b1110001110110,
13'b1110010000010,
13'b1110010000011,
13'b1110010000100,
13'b1110010000101,
13'b1110010000110,
13'b1110010010001,
13'b1110010010010,
13'b1110010010011,
13'b1110010010100,
13'b1110010010101,
13'b1110010010110,
13'b1110010100001,
13'b1110010100010,
13'b1110010100011,
13'b1110010100100,
13'b1110010100101,
13'b1110010100110,
13'b1110010110001,
13'b1110010110010,
13'b1110010110011,
13'b1110010110100,
13'b1110010110101,
13'b1110011000011,
13'b1110011000100,
13'b1111001110100,
13'b1111001110101,
13'b1111010000010,
13'b1111010000011,
13'b1111010000100,
13'b1111010000101,
13'b1111010000110,
13'b1111010010001,
13'b1111010010010,
13'b1111010010011,
13'b1111010010100,
13'b1111010010101,
13'b1111010010110,
13'b1111010100001,
13'b1111010100010,
13'b1111010100011,
13'b1111010100100,
13'b1111010100101,
13'b1111010100110,
13'b1111010110001,
13'b1111010110010,
13'b1111010110011,
13'b1111010110100,
13'b1111010110101: edge_mask_reg_512p3[183] <= 1'b1;
 		default: edge_mask_reg_512p3[183] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10110010110,
13'b10110010111,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101110100110,
13'b101110100111,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001111000011,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1010111000011,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111110001,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111110001,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1100111010010,
13'b1100111010011,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111110001,
13'b1100111110010,
13'b1100111110011,
13'b1101111010010,
13'b1101111100001,
13'b1101111100010,
13'b1101111100011,
13'b1101111110001,
13'b1101111110010,
13'b1101111110011,
13'b1110111010010,
13'b1110111100000,
13'b1110111100001,
13'b1110111100010,
13'b1110111110000,
13'b1110111110001,
13'b1110111110010,
13'b1111111010001,
13'b1111111010010,
13'b1111111100001,
13'b1111111100010,
13'b1111111110000,
13'b1111111110001,
13'b1111111110010: edge_mask_reg_512p3[184] <= 1'b1;
 		default: edge_mask_reg_512p3[184] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101101000,
13'b10101101001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101111000,
13'b101101111001,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110001000,
13'b110110001001,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111101000,
13'b1000110010011,
13'b1000110010100,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1001110100011,
13'b1001110100100,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1010110110011,
13'b1010110110100,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111100001,
13'b1010111100011: edge_mask_reg_512p3[185] <= 1'b1;
 		default: edge_mask_reg_512p3[185] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110101,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b100001100101,
13'b100001100110,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b101001100110,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110110,
13'b101100110111,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110110,
13'b110100110111,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100010011,
13'b111100010100,
13'b1000010010010,
13'b1000010010011,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1001010010001,
13'b1001010010010,
13'b1001010010011,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010110000,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1010010010001,
13'b1010010010010,
13'b1010010010011,
13'b1010010100000,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010110000,
13'b1010010110001,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010011000000,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100010001,
13'b1010100010010,
13'b1011010010001,
13'b1011010010010,
13'b1011010100000,
13'b1011010100001,
13'b1011010100010,
13'b1011010100011,
13'b1011010110000,
13'b1011010110001,
13'b1011010110010,
13'b1011010110011,
13'b1011011000000,
13'b1011011000001,
13'b1011011000010,
13'b1011011000011,
13'b1011011010000,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1100010010001,
13'b1100010010010,
13'b1100010100000,
13'b1100010100001,
13'b1100010100010,
13'b1100010110000,
13'b1100010110001,
13'b1100010110010,
13'b1100011000000,
13'b1100011000001,
13'b1100011000010,
13'b1100011000011,
13'b1100011010000,
13'b1100011010001,
13'b1100011010010,
13'b1100011010011,
13'b1100011100000,
13'b1100011100001,
13'b1100011100010,
13'b1100011100011,
13'b1100011110000,
13'b1100011110001,
13'b1100011110010,
13'b1100100000000,
13'b1100100000001,
13'b1101010100000,
13'b1101010100001,
13'b1101010110000,
13'b1101010110001,
13'b1101011000000,
13'b1101011000001,
13'b1101011010000,
13'b1101011010001,
13'b1101011100000,
13'b1101011100001,
13'b1101011110000,
13'b1101011110001,
13'b1110010100000,
13'b1110010110000,
13'b1110011000000,
13'b1110011010000,
13'b1110011100000,
13'b1110011110000: edge_mask_reg_512p3[186] <= 1'b1;
 		default: edge_mask_reg_512p3[186] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001101011,
13'b1001101100,
13'b1001111011,
13'b1001111100,
13'b10001011011,
13'b10001011100,
13'b10001101011,
13'b10001101100,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000: edge_mask_reg_512p3[187] <= 1'b1;
 		default: edge_mask_reg_512p3[187] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010111,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010110,
13'b100001010111,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000110,
13'b110001000111,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000100110,
13'b111000100111,
13'b1000000010110,
13'b1000000010111,
13'b1000000011000,
13'b1001000010110,
13'b1001000010111,
13'b1001000011000,
13'b1010000000110,
13'b1010000000111,
13'b1010000001000,
13'b1010000010110,
13'b1010000010111,
13'b1010000011000,
13'b1010000100110,
13'b1010000100111,
13'b1011000000110,
13'b1011000000111,
13'b1011000001000,
13'b1011000010110,
13'b1011000010111,
13'b1011000011000,
13'b1011000100110,
13'b1011000100111,
13'b1100000000110,
13'b1100000000111,
13'b1100000001000,
13'b1100000010110,
13'b1100000010111,
13'b1100000011000,
13'b1100000100111,
13'b1101000000100,
13'b1101000000101,
13'b1101000000110,
13'b1101000000111,
13'b1101000001000,
13'b1101000010100,
13'b1101000010101,
13'b1101000010110,
13'b1101000010111,
13'b1101000011000,
13'b1101000100110,
13'b1101000100111,
13'b1110000000100,
13'b1110000000101,
13'b1110000000110,
13'b1110000000111,
13'b1110000001000,
13'b1110000010100,
13'b1110000010101,
13'b1110000010110,
13'b1110000010111,
13'b1110000011000,
13'b1110000100110,
13'b1111000000100,
13'b1111000000101,
13'b1111000000110,
13'b1111000000111,
13'b1111000001000,
13'b1111000010100,
13'b1111000010101,
13'b1111000010110,
13'b1111000010111,
13'b1111000011000,
13'b1111000100110: edge_mask_reg_512p3[188] <= 1'b1;
 		default: edge_mask_reg_512p3[188] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b100010111010,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b101011001001,
13'b101011001010,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b110011101001,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110001001,
13'b110110011001,
13'b111011111000,
13'b111011111001,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b1000011101000,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101110111,
13'b1000101111000,
13'b1001011101000,
13'b1001011110111,
13'b1001011111000,
13'b1001011111001,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100010111,
13'b1001100011000,
13'b1001100011001,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1010011101000,
13'b1010011110111,
13'b1010011111000,
13'b1010011111001,
13'b1010100000111,
13'b1010100001000,
13'b1010100001001,
13'b1010100010111,
13'b1010100011000,
13'b1010100011001,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100101001,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1011011110111,
13'b1011011111000,
13'b1011011111001,
13'b1011100000110,
13'b1011100000111,
13'b1011100001000,
13'b1011100001001,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100011001,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100101001,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1100011110111,
13'b1100011111000,
13'b1100100000110,
13'b1100100000111,
13'b1100100001000,
13'b1100100001001,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1100100011001,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100101,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1101011110111,
13'b1101011111000,
13'b1101011111001,
13'b1101100000111,
13'b1101100001000,
13'b1101100001001,
13'b1101100010110,
13'b1101100010111,
13'b1101100011000,
13'b1101100011001,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100101001,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101100111001,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110110,
13'b1101101110111,
13'b1110011111000,
13'b1110011111001,
13'b1110100000111,
13'b1110100001000,
13'b1110100001001,
13'b1110100010111,
13'b1110100011000,
13'b1110100011001,
13'b1110100100111,
13'b1110100101000,
13'b1110100101001,
13'b1110100110110,
13'b1110100110111,
13'b1110100111000,
13'b1110100111001,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101001001,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110110,
13'b1110101110111,
13'b1111011111001,
13'b1111100000111,
13'b1111100001000,
13'b1111100001001,
13'b1111100001010,
13'b1111100010111,
13'b1111100011000,
13'b1111100011001,
13'b1111100011010,
13'b1111100100111,
13'b1111100101000,
13'b1111100101001,
13'b1111100110111,
13'b1111100111000,
13'b1111100111001,
13'b1111101000110,
13'b1111101000111,
13'b1111101001000,
13'b1111101001001,
13'b1111101010110,
13'b1111101010111,
13'b1111101011000,
13'b1111101011001,
13'b1111101100110,
13'b1111101100111,
13'b1111101101000: edge_mask_reg_512p3[189] <= 1'b1;
 		default: edge_mask_reg_512p3[189] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101101101001,
13'b101101101010,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001001,
13'b101111001010,
13'b101111011001,
13'b101111011010,
13'b110110001001,
13'b110110001010,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b110111001001,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110111001,
13'b111110111010,
13'b1000110001001,
13'b1000110001010,
13'b1000110001011,
13'b1000110011001,
13'b1000110011010,
13'b1000110011011,
13'b1000110101000,
13'b1000110101001,
13'b1000110101010,
13'b1000110111000,
13'b1000110111001,
13'b1000110111010,
13'b1000111001010,
13'b1001110001001,
13'b1001110001010,
13'b1001110001011,
13'b1001110011001,
13'b1001110011010,
13'b1001110011011,
13'b1001110101000,
13'b1001110101001,
13'b1001110101010,
13'b1001110111000,
13'b1001110111001,
13'b1001110111010,
13'b1001111001001,
13'b1001111001010,
13'b1010110001001,
13'b1010110001010,
13'b1010110001011,
13'b1010110011001,
13'b1010110011010,
13'b1010110011011,
13'b1010110101000,
13'b1010110101001,
13'b1010110101010,
13'b1010110111000,
13'b1010110111001,
13'b1010110111010,
13'b1010111001010,
13'b1011110001001,
13'b1011110001010,
13'b1011110001011,
13'b1011110011001,
13'b1011110011010,
13'b1011110011011,
13'b1011110101000,
13'b1011110101001,
13'b1011110101010,
13'b1011110111000,
13'b1011110111001,
13'b1011110111010,
13'b1100110001001,
13'b1100110001010,
13'b1100110001011,
13'b1100110011000,
13'b1100110011001,
13'b1100110011010,
13'b1100110011011,
13'b1100110101000,
13'b1100110101001,
13'b1100110101010,
13'b1100110101011,
13'b1100110111000,
13'b1100110111001,
13'b1100110111010,
13'b1100111001001,
13'b1101110001001,
13'b1101110001010,
13'b1101110001011,
13'b1101110011000,
13'b1101110011001,
13'b1101110011010,
13'b1101110011011,
13'b1101110101000,
13'b1101110101001,
13'b1101110101010,
13'b1101110101011,
13'b1101110111000,
13'b1101110111001,
13'b1101110111010,
13'b1101111001001,
13'b1110110001001,
13'b1110110001010,
13'b1110110011000,
13'b1110110011001,
13'b1110110011010,
13'b1110110101000,
13'b1110110101001,
13'b1110110101010,
13'b1110110111000,
13'b1110110111001,
13'b1110110111010,
13'b1111110011000,
13'b1111110011001,
13'b1111110011010,
13'b1111110101000,
13'b1111110101001,
13'b1111110101010: edge_mask_reg_512p3[190] <= 1'b1;
 		default: edge_mask_reg_512p3[190] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[191] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[192] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b11001000000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100111,
13'b11010101000,
13'b100000110000,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000000,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010000,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100111,
13'b100010101000,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100000,
13'b101001100001,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100111,
13'b101010101000,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110000,
13'b110001110001,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010111,
13'b110010011000,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010110,
13'b111000010111,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1010000110010,
13'b1010000110011,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010010,
13'b1010001010011,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1011001010011,
13'b1011001100010,
13'b1011001100011,
13'b1011001110011: edge_mask_reg_512p3[193] <= 1'b1;
 		default: edge_mask_reg_512p3[193] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b11001000000,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010000,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000101,
13'b11011000110,
13'b100000110000,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000000,
13'b100001000001,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010000,
13'b100001010001,
13'b100001010010,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100000,
13'b100001100001,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110000,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000000,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100011000101,
13'b100011000110,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101011000101,
13'b101011000110,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100000,
13'b110010100001,
13'b110010100101,
13'b110010100110,
13'b110010110101,
13'b110010110110,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010110,
13'b111000010111,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100110,
13'b111000100111,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110110,
13'b111000110111,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000110,
13'b111001000111,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000101,
13'b111010000110,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010100001,
13'b1000000010000,
13'b1000000010001,
13'b1000000100000,
13'b1000000100001,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001110000,
13'b1000001110001,
13'b1000010000000,
13'b1000010000001,
13'b1000010010000,
13'b1000010010001: edge_mask_reg_512p3[194] <= 1'b1;
 		default: edge_mask_reg_512p3[194] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101001001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111001,
13'b10100111010,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b101001001001,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b101100011010,
13'b110001100110,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b111001100110,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1001001100100,
13'b1001001100101,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1011001110100,
13'b1011001110101,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010010110,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010110011,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110110,
13'b1101010000011,
13'b1101010000100,
13'b1101010010011,
13'b1101010010100,
13'b1101010010101,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010110011,
13'b1101010110100,
13'b1101010110101,
13'b1101010110110,
13'b1101011000011,
13'b1101011000100,
13'b1101011000101,
13'b1101011000110,
13'b1101011010100,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011100101,
13'b1101011100110,
13'b1101011100111,
13'b1110010010100,
13'b1110010100100,
13'b1110010100101,
13'b1110010110100,
13'b1110010110101,
13'b1110010110110,
13'b1110011000100,
13'b1110011000101,
13'b1110011000110,
13'b1110011010100,
13'b1110011010101,
13'b1110011010110,
13'b1110011010111,
13'b1110011100100,
13'b1110011100101,
13'b1110011100110,
13'b1111010110101,
13'b1111011000101,
13'b1111011000110,
13'b1111011010101,
13'b1111011010110,
13'b1111011100101,
13'b1111011100110: edge_mask_reg_512p3[195] <= 1'b1;
 		default: edge_mask_reg_512p3[195] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11011100,
13'b11101011,
13'b11101100,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b11111101,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100001101,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100011101,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100101101,
13'b100111010,
13'b100111011,
13'b100111100,
13'b100111101,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101001101,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101011101,
13'b101101010,
13'b101101011,
13'b101101100,
13'b101101101,
13'b1011111011,
13'b1011111100,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100001101,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100011101,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100101101,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101001101,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101011101,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101101101,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1101111101,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110001101,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b1110011101,
13'b10100011011,
13'b10100011100,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11100111001,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111010,
13'b11110111011,
13'b100100111000,
13'b100100111001,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100101111100,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111010,
13'b100110111011,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111010,
13'b101110111011,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111010,
13'b111101000111,
13'b111101001000,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110111010,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1000110001010,
13'b1000110001011,
13'b1000110011000,
13'b1000110011001,
13'b1000110011010,
13'b1000110011011,
13'b1000110101001,
13'b1000110101010,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001101111001,
13'b1001101111010,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110001001,
13'b1001110001010,
13'b1001110010111,
13'b1001110011000,
13'b1001110011001,
13'b1001110011010,
13'b1010101010110,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010101111001,
13'b1010101111010,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110001001,
13'b1010110001010,
13'b1010110010111,
13'b1010110011000,
13'b1010110011001,
13'b1010110011010,
13'b1011101100111,
13'b1011101101000,
13'b1011101110111,
13'b1011101111000,
13'b1011101111001,
13'b1011110000111,
13'b1011110001000,
13'b1011110001001,
13'b1011110001010,
13'b1011110011000,
13'b1011110011001,
13'b1011110011010: edge_mask_reg_512p3[196] <= 1'b1;
 		default: edge_mask_reg_512p3[196] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110000,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110010,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101101000110,
13'b101101000111,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111010000,
13'b1000101100010,
13'b1000101100011,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000111000000,
13'b1000111000001,
13'b1001101100011,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110110001,
13'b1010110110010,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1100110000000,
13'b1100110000001,
13'b1100110010000: edge_mask_reg_512p3[197] <= 1'b1;
 		default: edge_mask_reg_512p3[197] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000101,
13'b100010000110,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000101,
13'b101010000110,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110101,
13'b110001110110,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010011,
13'b1000001010100,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000000101,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000000100,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000010100,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100000110100,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1100001000011,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000000100,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1101000010011,
13'b1101000010100,
13'b1101000100000,
13'b1101000100001,
13'b1101000100010,
13'b1101000100011,
13'b1101000110000,
13'b1101000110001,
13'b1101000110010,
13'b1101000110011,
13'b1101001000000,
13'b1101001000001,
13'b1101001000010,
13'b1101001000011,
13'b1101001010000,
13'b1101001010001,
13'b1101001010010,
13'b1101001010011,
13'b1110000000000,
13'b1110000000001,
13'b1110000000010,
13'b1110000000011,
13'b1110000010000,
13'b1110000010001,
13'b1110000010010,
13'b1110000010011,
13'b1110000100000,
13'b1110000100001,
13'b1110000100010,
13'b1110000100011,
13'b1110000110000,
13'b1110000110001,
13'b1110000110010,
13'b1110000110011,
13'b1110001000000,
13'b1110001000001,
13'b1110001000010,
13'b1110001010000,
13'b1111000000000,
13'b1111000000001,
13'b1111000000010,
13'b1111000010000,
13'b1111000010001,
13'b1111000010010,
13'b1111000100000,
13'b1111000100001,
13'b1111000100010,
13'b1111000110000,
13'b1111000110001,
13'b1111001000000,
13'b1111001000001: edge_mask_reg_512p3[198] <= 1'b1;
 		default: edge_mask_reg_512p3[198] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000101,
13'b100010000110,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000101,
13'b101010000110,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001100101,
13'b110001100110,
13'b110001110101,
13'b110001110110,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1100001000011,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1101000100000,
13'b1101000100001,
13'b1101000100010,
13'b1101000100011,
13'b1101000110000,
13'b1101000110001,
13'b1101000110010,
13'b1101000110011,
13'b1101001000000,
13'b1101001000001,
13'b1101001000010,
13'b1101001000011,
13'b1101001010000,
13'b1101001010001,
13'b1101001010010,
13'b1101001010011,
13'b1110000000000,
13'b1110000000001,
13'b1110000010000,
13'b1110000010001,
13'b1110000100000,
13'b1110000100001,
13'b1110000110000,
13'b1110000110001,
13'b1110000110010,
13'b1110001000000,
13'b1110001000001,
13'b1110001000010,
13'b1110001010000,
13'b1111000010000,
13'b1111000100000,
13'b1111000110000,
13'b1111000110001,
13'b1111001000000,
13'b1111001000001: edge_mask_reg_512p3[199] <= 1'b1;
 		default: edge_mask_reg_512p3[199] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010111,
13'b1010011000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b11001000000,
13'b11001000001,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010000,
13'b11001010001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100000,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b100000110000,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000000,
13'b100001000001,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010000,
13'b100001010001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100000,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000111,
13'b100010001000,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100000,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000111,
13'b101010001000,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100000,
13'b110001100001,
13'b110001100011,
13'b110001100100,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110111,
13'b110001111000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010111,
13'b111000011000,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100111,
13'b111000101000,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001100010,
13'b111001100011,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001100010,
13'b1000001100011,
13'b1001000100010,
13'b1001000100011,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001010010,
13'b1001001010011: edge_mask_reg_512p3[200] <= 1'b1;
 		default: edge_mask_reg_512p3[200] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100001000,
13'b1100001001,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100111,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010111,
13'b110101011000,
13'b111011100110,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110100,
13'b111100110101,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110011,
13'b1001100110100,
13'b1010011100011,
13'b1010011100100,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1011011100011,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1100011110001,
13'b1100011110010,
13'b1100011110011,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100000100,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1101011110001,
13'b1101011110010,
13'b1101100000000,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100100001,
13'b1101100100010,
13'b1110011110001,
13'b1110100000001,
13'b1110100000010,
13'b1110100010001,
13'b1110100010010,
13'b1110100100001,
13'b1111100010001,
13'b1111100010010: edge_mask_reg_512p3[201] <= 1'b1;
 		default: edge_mask_reg_512p3[201] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110101,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110101,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100111,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000010,
13'b110011000011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010111,
13'b111011000010,
13'b111011000011,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011100000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110100,
13'b111100110101,
13'b1000011000001,
13'b1000011000010,
13'b1000011010000,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110011,
13'b1001100110100,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1011011010001,
13'b1011011010010,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1100011100000,
13'b1100011100001,
13'b1100011110000,
13'b1100011110001,
13'b1100011110010,
13'b1100011110011,
13'b1100100000000,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100010000,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1101011100000,
13'b1101011110000,
13'b1101011110001,
13'b1101011110010,
13'b1101100000000,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100100001,
13'b1101100100010,
13'b1110011110000,
13'b1110011110001,
13'b1110100000000,
13'b1110100000001,
13'b1110100000010,
13'b1110100010000,
13'b1110100010001,
13'b1110100010010,
13'b1110100100001,
13'b1111100010001,
13'b1111100010010: edge_mask_reg_512p3[202] <= 1'b1;
 		default: edge_mask_reg_512p3[202] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b110011011000,
13'b110011011001,
13'b110011101000,
13'b110011101001,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011001,
13'b111011101001,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b1000011101010,
13'b1000011111000,
13'b1000011111001,
13'b1000011111010,
13'b1000100001000,
13'b1000100001001,
13'b1000100001010,
13'b1000100001011,
13'b1000100011000,
13'b1000100011001,
13'b1000100011010,
13'b1000100011011,
13'b1000100101001,
13'b1000100101010,
13'b1000100101011,
13'b1000100111001,
13'b1000100111010,
13'b1000100111011,
13'b1000101001011,
13'b1001011101010,
13'b1001011111000,
13'b1001011111001,
13'b1001011111010,
13'b1001011111011,
13'b1001100001000,
13'b1001100001001,
13'b1001100001010,
13'b1001100001011,
13'b1001100011001,
13'b1001100011010,
13'b1001100011011,
13'b1001100101001,
13'b1001100101010,
13'b1001100101011,
13'b1001100111001,
13'b1001100111010,
13'b1001100111011,
13'b1001101001011,
13'b1010011101010,
13'b1010011111001,
13'b1010011111010,
13'b1010011111011,
13'b1010100001001,
13'b1010100001010,
13'b1010100001011,
13'b1010100001100,
13'b1010100011001,
13'b1010100011010,
13'b1010100011011,
13'b1010100011100,
13'b1010100101001,
13'b1010100101010,
13'b1010100101011,
13'b1010100101100,
13'b1010100111001,
13'b1010100111010,
13'b1010100111011,
13'b1010100111100,
13'b1010101001011,
13'b1011011101001,
13'b1011011101010,
13'b1011011111001,
13'b1011011111010,
13'b1011011111011,
13'b1011100001001,
13'b1011100001010,
13'b1011100001011,
13'b1011100001100,
13'b1011100011001,
13'b1011100011010,
13'b1011100011011,
13'b1011100011100,
13'b1011100101001,
13'b1011100101010,
13'b1011100101011,
13'b1011100101100,
13'b1011100111010,
13'b1011100111011,
13'b1011100111100,
13'b1011101001011,
13'b1011101001100,
13'b1100011101010,
13'b1100011111001,
13'b1100011111010,
13'b1100011111011,
13'b1100100001001,
13'b1100100001010,
13'b1100100001011,
13'b1100100001100,
13'b1100100011001,
13'b1100100011010,
13'b1100100011011,
13'b1100100011100,
13'b1100100101001,
13'b1100100101010,
13'b1100100101011,
13'b1100100101100,
13'b1100100111010,
13'b1100100111011,
13'b1100100111100,
13'b1100101001011,
13'b1100101001100,
13'b1101011101010,
13'b1101011111001,
13'b1101011111010,
13'b1101011111011,
13'b1101100001001,
13'b1101100001010,
13'b1101100001011,
13'b1101100001100,
13'b1101100011001,
13'b1101100011010,
13'b1101100011011,
13'b1101100011100,
13'b1101100101001,
13'b1101100101010,
13'b1101100101011,
13'b1101100101100,
13'b1101100101101,
13'b1101100111010,
13'b1101100111011,
13'b1101100111100,
13'b1110011111001,
13'b1110011111010,
13'b1110011111011,
13'b1110100001001,
13'b1110100001010,
13'b1110100001011,
13'b1110100001100,
13'b1110100011001,
13'b1110100011010,
13'b1110100011011,
13'b1110100011100,
13'b1110100011101,
13'b1110100101010,
13'b1110100101011,
13'b1110100101100,
13'b1110100101101,
13'b1110100111010,
13'b1110100111011,
13'b1110100111100,
13'b1110100111101,
13'b1111011111010,
13'b1111011111011,
13'b1111100001010,
13'b1111100001011,
13'b1111100001100,
13'b1111100011010,
13'b1111100011011,
13'b1111100011100,
13'b1111100011101,
13'b1111100101011,
13'b1111100101100,
13'b1111100101101,
13'b1111100111100,
13'b1111100111101: edge_mask_reg_512p3[203] <= 1'b1;
 		default: edge_mask_reg_512p3[203] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b110011001000,
13'b110011001001,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011101011,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110011111011,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b111011011001,
13'b111011011010,
13'b111011011011,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011101011,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111011111011,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100101001,
13'b1000011011001,
13'b1000011011010,
13'b1000011011011,
13'b1000011101001,
13'b1000011101010,
13'b1000011101011,
13'b1000011111000,
13'b1000011111001,
13'b1000011111010,
13'b1000011111011,
13'b1000100001000,
13'b1000100001001,
13'b1000100001010,
13'b1000100001011,
13'b1000100011000,
13'b1000100011001,
13'b1000100011010,
13'b1000100011011,
13'b1001011011001,
13'b1001011011010,
13'b1001011011011,
13'b1001011101001,
13'b1001011101010,
13'b1001011101011,
13'b1001011111000,
13'b1001011111001,
13'b1001011111010,
13'b1001011111011,
13'b1001100001000,
13'b1001100001001,
13'b1001100001010,
13'b1001100001011,
13'b1001100011001,
13'b1001100011010,
13'b1001100011011,
13'b1001100101001,
13'b1001100101010,
13'b1010011011001,
13'b1010011011010,
13'b1010011011011,
13'b1010011101001,
13'b1010011101010,
13'b1010011101011,
13'b1010011111001,
13'b1010011111010,
13'b1010011111011,
13'b1010100001001,
13'b1010100001010,
13'b1010100001011,
13'b1010100011001,
13'b1010100011010,
13'b1010100011011,
13'b1010100101001,
13'b1010100101010,
13'b1011011011010,
13'b1011011011011,
13'b1011011101001,
13'b1011011101010,
13'b1011011101011,
13'b1011011101100,
13'b1011011111001,
13'b1011011111010,
13'b1011011111011,
13'b1011011111100,
13'b1011100001001,
13'b1011100001010,
13'b1011100001011,
13'b1011100011001,
13'b1011100011010,
13'b1011100011011,
13'b1011100101001,
13'b1011100101010,
13'b1100011011010,
13'b1100011011011,
13'b1100011011100,
13'b1100011101001,
13'b1100011101010,
13'b1100011101011,
13'b1100011101100,
13'b1100011111001,
13'b1100011111010,
13'b1100011111011,
13'b1100011111100,
13'b1100100001001,
13'b1100100001010,
13'b1100100001011,
13'b1100100001100,
13'b1100100011001,
13'b1100100011010,
13'b1100100011011,
13'b1100100101010,
13'b1100100101011,
13'b1101011011010,
13'b1101011011011,
13'b1101011011100,
13'b1101011101001,
13'b1101011101010,
13'b1101011101011,
13'b1101011101100,
13'b1101011111001,
13'b1101011111010,
13'b1101011111011,
13'b1101011111100,
13'b1101100001001,
13'b1101100001010,
13'b1101100001011,
13'b1101100001100,
13'b1101100011001,
13'b1101100011010,
13'b1101100011011,
13'b1101100101001,
13'b1101100101010,
13'b1101100101011,
13'b1110011011010,
13'b1110011011011,
13'b1110011101001,
13'b1110011101010,
13'b1110011101011,
13'b1110011101100,
13'b1110011111001,
13'b1110011111010,
13'b1110011111011,
13'b1110011111100,
13'b1110100001001,
13'b1110100001010,
13'b1110100001011,
13'b1110100001100,
13'b1110100011001,
13'b1110100011010,
13'b1110100011011,
13'b1110100101010,
13'b1111011101010,
13'b1111011101011,
13'b1111011101100,
13'b1111011111010,
13'b1111011111011,
13'b1111011111100,
13'b1111100001010,
13'b1111100001011,
13'b1111100001100,
13'b1111100011010,
13'b1111100011011: edge_mask_reg_512p3[204] <= 1'b1;
 		default: edge_mask_reg_512p3[204] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[205] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010100,
13'b10010101,
13'b10010110,
13'b10100100,
13'b10100101,
13'b10100110,
13'b10110101,
13'b10110110,
13'b11000100,
13'b11000101,
13'b11000110,
13'b11010100,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100100,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110100,
13'b11110101,
13'b11110110,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100010100,
13'b100010101,
13'b100010110,
13'b100100100,
13'b100100101,
13'b100100110,
13'b100110100,
13'b100110101,
13'b100110110,
13'b1001100100,
13'b1001100101,
13'b1001100110,
13'b1001110100,
13'b1001110101,
13'b1001110110,
13'b1010000100,
13'b1010000101,
13'b1010000110,
13'b1010010100,
13'b1010010101,
13'b1010010110,
13'b1010100100,
13'b1010100101,
13'b1010100110,
13'b1010110100,
13'b1010110101,
13'b1010110110,
13'b1011000011,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011010011,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011100011,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100110100,
13'b1100110101,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001100011,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001110011,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10010000011,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010010011,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010100011,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010110011,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10011000010,
13'b10011000011,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011010010,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011100010,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b11001000011,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010010001,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010100000,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010110000,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11011000000,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011010000,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011100000,
13'b11011100001,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011110000,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11100000000,
13'b11100000001,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100010000000,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010010000,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010100000,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010110000,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100011000000,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011110000,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100100000000,
13'b100100000001,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100100,
13'b100100100101,
13'b101001000100,
13'b101001000101,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101011000000,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011110000,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101100000000,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100100100,
13'b101100100101,
13'b110001010100,
13'b110001010101,
13'b110001100000,
13'b110001100100,
13'b110001100101,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110011000000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011010000,
13'b110011010001,
13'b110011010010,
13'b110011010100,
13'b110011010101,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100100,
13'b110011100101,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110100,
13'b110011110101,
13'b110100000100,
13'b110100000101,
13'b111001100000,
13'b111001100001,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111011000000,
13'b111011000001,
13'b111011000010,
13'b111011010000,
13'b111011010001,
13'b111011100000,
13'b111011100001,
13'b1000001100000,
13'b1000001110000,
13'b1000001110001,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010010000,
13'b1000010010001,
13'b1000010010010,
13'b1000010100000,
13'b1000010100001,
13'b1000010100010,
13'b1000010110000,
13'b1000010110001,
13'b1000010110010,
13'b1000011000000,
13'b1000011000001,
13'b1000011010000,
13'b1001001100000,
13'b1001001110000,
13'b1001010000000,
13'b1001010010000,
13'b1001010010001,
13'b1001010100000,
13'b1001010100001,
13'b1001010110000,
13'b1001011000000,
13'b1010010000000,
13'b1010010010000,
13'b1010010100000,
13'b1010010110000: edge_mask_reg_512p3[206] <= 1'b1;
 		default: edge_mask_reg_512p3[206] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000100101,
13'b101000100110: edge_mask_reg_512p3[207] <= 1'b1;
 		default: edge_mask_reg_512p3[207] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[208] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100001000,
13'b100100001001,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001001,
13'b101111001010,
13'b110100011000,
13'b110100011001,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010111,
13'b111110011000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110010110,
13'b1000110010111,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010110,
13'b1001110010111,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1011100110101,
13'b1011100110110,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011101110111,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1100100110101,
13'b1100100110110,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101100110,
13'b1100101100111,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100101110110,
13'b1100101110111,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110000111,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1101101000100,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101010011,
13'b1101101010100,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101100011,
13'b1101101100100,
13'b1101101100101,
13'b1101101100110,
13'b1101101100111,
13'b1101101110011,
13'b1101101110100,
13'b1101101110101,
13'b1101101110110,
13'b1101101110111,
13'b1101110000011,
13'b1101110000100,
13'b1101110000101,
13'b1101110000110,
13'b1101110000111,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1101110010110,
13'b1110101010011,
13'b1110101010100,
13'b1110101010101,
13'b1110101010110,
13'b1110101100011,
13'b1110101100100,
13'b1110101100101,
13'b1110101110011,
13'b1110101110100,
13'b1110101110101,
13'b1110110000011,
13'b1110110000100,
13'b1110110000101,
13'b1110110010100,
13'b1110110010101,
13'b1111101010100,
13'b1111101010101,
13'b1111101100100,
13'b1111101100101,
13'b1111101110100: edge_mask_reg_512p3[209] <= 1'b1;
 		default: edge_mask_reg_512p3[209] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11100101001,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100100101001,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101100111001,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011001,
13'b101111011010,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111001000,
13'b110111001001,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000111,
13'b111111001000,
13'b1000101010111,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110011001,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000111000111,
13'b1000111001000,
13'b1001101010111,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001110111001,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010110111000,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011101110111,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011110111000,
13'b1011111000110,
13'b1011111000111,
13'b1100101100101,
13'b1100101100110,
13'b1100101110100,
13'b1100101110101,
13'b1100101110110,
13'b1100101110111,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110000111,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1100110100100,
13'b1100110100101,
13'b1100110100110,
13'b1100110100111,
13'b1100110110100,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000100,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1101101110100,
13'b1101101110101,
13'b1101101110110,
13'b1101110000011,
13'b1101110000100,
13'b1101110000101,
13'b1101110000110,
13'b1101110000111,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1101110010110,
13'b1101110010111,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1101110110100,
13'b1101110110101,
13'b1101110110110,
13'b1101111000100,
13'b1101111000101,
13'b1110101110100,
13'b1110110000011,
13'b1110110000100,
13'b1110110010100,
13'b1110110010101,
13'b1110110100100,
13'b1110110100101,
13'b1110110110100,
13'b1110110110101: edge_mask_reg_512p3[210] <= 1'b1;
 		default: edge_mask_reg_512p3[210] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11100101001,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100100101001,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101100111001,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011001,
13'b101111011010,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110111000,
13'b110110111001,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110111000,
13'b1000101010111,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110011001,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110110111,
13'b1000110111000,
13'b1001101010111,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110011001,
13'b1001110100111,
13'b1001110101000,
13'b1001110101001,
13'b1001110110111,
13'b1001110111000,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110111,
13'b1010110111000,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011101110111,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110110110,
13'b1011110110111,
13'b1100101100101,
13'b1100101100110,
13'b1100101110100,
13'b1100101110101,
13'b1100101110110,
13'b1100101110111,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110000111,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1100110100101,
13'b1100110100110,
13'b1100110100111,
13'b1100110101000,
13'b1100110110110,
13'b1100110110111,
13'b1101101110100,
13'b1101101110101,
13'b1101101110110,
13'b1101110000011,
13'b1101110000100,
13'b1101110000101,
13'b1101110000110,
13'b1101110000111,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1101110010110,
13'b1101110010111,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1101110100111,
13'b1101110101000,
13'b1101110110111,
13'b1110101110100,
13'b1110101110101,
13'b1110110000011,
13'b1110110000100,
13'b1110110000101,
13'b1110110000110,
13'b1110110010100,
13'b1110110010101,
13'b1110110010110,
13'b1110110100100,
13'b1110110100101,
13'b1110110100110,
13'b1111110000100,
13'b1111110000101,
13'b1111110010100,
13'b1111110010101,
13'b1111110010110,
13'b1111110100101,
13'b1111110100110: edge_mask_reg_512p3[211] <= 1'b1;
 		default: edge_mask_reg_512p3[211] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b1010000000010: edge_mask_reg_512p3[212] <= 1'b1;
 		default: edge_mask_reg_512p3[212] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110111,
13'b100111000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011100110,
13'b1011100111,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100000,
13'b11011100001,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110000,
13'b11011110001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000000,
13'b11100000001,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100101000,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100011,
13'b100010100100,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110000,
13'b100011110001,
13'b100011110010,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000000,
13'b100100000001,
13'b100100000010,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010000,
13'b100100010001,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b101010000111,
13'b101010001000,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110000,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000000,
13'b101100000001,
13'b101100000010,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010000,
13'b101100010001,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100001,
13'b110010100010,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010000,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010000,
13'b110100010001,
13'b110100010111,
13'b110100011000,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010000,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111100000000,
13'b111100000001,
13'b1000010110010,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011100001,
13'b1001011100010: edge_mask_reg_512p3[213] <= 1'b1;
 		default: edge_mask_reg_512p3[213] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[214] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[215] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[216] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[217] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[218] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010100,
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100100,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010100,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100100,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010100,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100100,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1001100100,
13'b1001100101,
13'b1001100110,
13'b1001110100,
13'b1001110101,
13'b1001110110,
13'b1010000100,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010100,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100100,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110100,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b10001010011,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001100011,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001110000,
13'b10001110001,
13'b10001110011,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10010000000,
13'b10010000001,
13'b10010000010,
13'b10010000011,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010010000,
13'b10010010001,
13'b10010010010,
13'b10010010011,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010100000,
13'b10010100001,
13'b10010100010,
13'b10010100011,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110000,
13'b10010110001,
13'b10010110010,
13'b10010110011,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000000,
13'b10011000001,
13'b10011000010,
13'b10011000011,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010001,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001110000,
13'b11001110001,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11010000000,
13'b11010000001,
13'b11010000010,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010010000,
13'b11010010001,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010100000,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110000,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000000,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011010000,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011100000,
13'b11011100001,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010101,
13'b11101010110,
13'b100001010100,
13'b100001010101,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001110000,
13'b100001110001,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100010000000,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010010000,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010100000,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010110000,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100011000000,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110000,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000001,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010101,
13'b100101010110,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001110000,
13'b101001110001,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101011000000,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110000,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000000,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101010101,
13'b101101010110,
13'b110001110100,
13'b110001110101,
13'b110010000100,
13'b110010000101,
13'b110010010000,
13'b110010010001,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110011000000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011010000,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000101,
13'b110101000110,
13'b111010100000,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111010110100,
13'b111011000000,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011010000,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011100000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100101,
13'b111011100110,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b1000010110000,
13'b1000011000000,
13'b1000011000001,
13'b1000011010000,
13'b1000011010001,
13'b1000011010010,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1001011010000,
13'b1001011010001,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001100000000,
13'b1001100000001,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1010011100000,
13'b1010011100001,
13'b1010011110000,
13'b1010011110001,
13'b1010100000000,
13'b1010100000001,
13'b1010100010000,
13'b1010100010001,
13'b1010100100000,
13'b1010100100001,
13'b1011100000000: edge_mask_reg_512p3[219] <= 1'b1;
 		default: edge_mask_reg_512p3[219] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110000,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101101100101,
13'b101101100110,
13'b101101110000,
13'b101101110001,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111110000000,
13'b111110010000,
13'b111110010101,
13'b111110010110,
13'b111110100000,
13'b111110100001,
13'b111110100101,
13'b111110100110,
13'b111110110000,
13'b111110110001,
13'b111110110101,
13'b111110110110,
13'b111111000000,
13'b111111000001,
13'b111111000101,
13'b111111000110,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010101,
13'b111111010110,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100101,
13'b111111100110: edge_mask_reg_512p3[220] <= 1'b1;
 		default: edge_mask_reg_512p3[220] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[221] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100110,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100101,
13'b100110100110,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000010,
13'b110011000011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010101,
13'b110110010110,
13'b111011000010,
13'b111011000011,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011100000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010110,
13'b111101010111,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100110,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b1000011000001,
13'b1000011000010,
13'b1000011010000,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101110000,
13'b1001101110001,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100110000,
13'b1010100110001,
13'b1010101000000,
13'b1010101000001,
13'b1010101010000,
13'b1010101010001,
13'b1010101100000,
13'b1011011100000,
13'b1011011100001,
13'b1011011110000,
13'b1011011110001,
13'b1011100000000,
13'b1011100000001,
13'b1011100010000,
13'b1011100100000,
13'b1011100110000,
13'b1011101000000,
13'b1011101010000,
13'b1100011100000,
13'b1100011110000,
13'b1100100000000,
13'b1100100010000,
13'b1100100100000: edge_mask_reg_512p3[222] <= 1'b1;
 		default: edge_mask_reg_512p3[222] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111100,
13'b101001011,
13'b101001100,
13'b101011011,
13'b101011100,
13'b101011101,
13'b101101010,
13'b101101011,
13'b101101100,
13'b101101101,
13'b1110011001,
13'b1110011010,
13'b10110011001,
13'b10110011010,
13'b10110101001,
13'b10110101010,
13'b11110011001,
13'b11110101000,
13'b11110101001,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110100101,
13'b110110100110,
13'b110110101000,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000111000110,
13'b1000111000111,
13'b1000111010110,
13'b1000111010111,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000: edge_mask_reg_512p3[223] <= 1'b1;
 		default: edge_mask_reg_512p3[223] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001101101,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1001111101,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010001101,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001101101,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10001111101,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010001101,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b11001001010,
13'b11001001011,
13'b11001001100,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001010,
13'b11011001011,
13'b100001001010,
13'b100001001011,
13'b100001011010,
13'b100001011011,
13'b100001101010,
13'b100001101011,
13'b100001111010,
13'b100001111011,
13'b100010001010,
13'b100010001011,
13'b100010011010,
13'b100010011011,
13'b101001001010,
13'b101001001011,
13'b101001011010,
13'b101001011011,
13'b101001101010,
13'b101001101011,
13'b101001111010,
13'b101001111011,
13'b101010001010,
13'b101010001011,
13'b101010011010,
13'b101010011011,
13'b110001001010,
13'b110001011010,
13'b110001011011,
13'b110001011100,
13'b110001101010,
13'b110001101011,
13'b110001111001,
13'b110001111010,
13'b110001111011,
13'b110010001001,
13'b110010001010,
13'b110010001011,
13'b110010011001,
13'b110010011010,
13'b110010011011,
13'b111001001010,
13'b111001001011,
13'b111001011001,
13'b111001011010,
13'b111001011011,
13'b111001011100,
13'b111001101001,
13'b111001101010,
13'b111001101011,
13'b111001111001,
13'b111001111010,
13'b111001111011,
13'b111010001001,
13'b111010001010,
13'b111010001011,
13'b111010011001,
13'b111010011010,
13'b111010011011,
13'b1000001001010,
13'b1000001001011,
13'b1000001011001,
13'b1000001011010,
13'b1000001011011,
13'b1000001011100,
13'b1000001101001,
13'b1000001101010,
13'b1000001101011,
13'b1000001111001,
13'b1000001111010,
13'b1000001111011,
13'b1000010001001,
13'b1000010001010,
13'b1000010001011,
13'b1000010011001,
13'b1000010011010,
13'b1000010011011,
13'b1001001001010,
13'b1001001001011,
13'b1001001011001,
13'b1001001011010,
13'b1001001011011,
13'b1001001101001,
13'b1001001101010,
13'b1001001101011,
13'b1001001111001,
13'b1001001111010,
13'b1001001111011,
13'b1001010001001,
13'b1001010001010,
13'b1001010001011,
13'b1001010011001,
13'b1001010011010,
13'b1001010011011,
13'b1010001001010,
13'b1010001001011,
13'b1010001011001,
13'b1010001011010,
13'b1010001011011,
13'b1010001011100,
13'b1010001101001,
13'b1010001101010,
13'b1010001101011,
13'b1010001101100,
13'b1010001111001,
13'b1010001111010,
13'b1010001111011,
13'b1010010001001,
13'b1010010001010,
13'b1010010001011,
13'b1010010011001,
13'b1010010011010,
13'b1010010011011,
13'b1011001001010,
13'b1011001001011,
13'b1011001011001,
13'b1011001011010,
13'b1011001011011,
13'b1011001011100,
13'b1011001101000,
13'b1011001101001,
13'b1011001101010,
13'b1011001101011,
13'b1011001101100,
13'b1011001111000,
13'b1011001111001,
13'b1011001111010,
13'b1011001111011,
13'b1011010001001,
13'b1011010001010,
13'b1011010001011,
13'b1011010011001,
13'b1011010011010,
13'b1011010011011,
13'b1100001001010,
13'b1100001001011,
13'b1100001011001,
13'b1100001011010,
13'b1100001011011,
13'b1100001101000,
13'b1100001101001,
13'b1100001101010,
13'b1100001101011,
13'b1100001111000,
13'b1100001111001,
13'b1100001111010,
13'b1100001111011,
13'b1100010001000,
13'b1100010001001,
13'b1100010001010,
13'b1100010001011,
13'b1100010011010,
13'b1101001011001,
13'b1101001011010,
13'b1101001011011,
13'b1101001101000,
13'b1101001101001,
13'b1101001101010,
13'b1101001101011,
13'b1101001111000,
13'b1101001111001,
13'b1101001111010,
13'b1101010001000,
13'b1101010001001,
13'b1110001011000,
13'b1110001011001,
13'b1110001011010,
13'b1110001101000,
13'b1110001101001,
13'b1110001101010,
13'b1110001111000,
13'b1110001111001,
13'b1110001111010,
13'b1110010001000,
13'b1110010001001,
13'b1111001011001,
13'b1111001011010,
13'b1111001101001,
13'b1111001101010,
13'b1111001111001,
13'b1111001111010: edge_mask_reg_512p3[224] <= 1'b1;
 		default: edge_mask_reg_512p3[224] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100111,
13'b1101110110,
13'b1101110111,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101100010110,
13'b101100010111,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000000,
13'b101110000001,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010000,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010000,
13'b110110010001,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100100,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b111100110001,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010111,
13'b111101011000,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100111,
13'b111101101000,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110100000,
13'b111110100001,
13'b111110100011,
13'b111110100100,
13'b1000101000001,
13'b1000101000010,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100000,
13'b1000110100010,
13'b1000110100011,
13'b1001101010001,
13'b1001101010010,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100010,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011: edge_mask_reg_512p3[225] <= 1'b1;
 		default: edge_mask_reg_512p3[225] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[226] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[227] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100111001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b10100101010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101001,
13'b11100101010,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110011,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110011,
13'b111011110100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110011,
13'b1000011110100,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011100101,
13'b1011011100110,
13'b1100010100101,
13'b1100010100110,
13'b1100010110101,
13'b1100010110110,
13'b1100011000101,
13'b1100011000110,
13'b1100011010101,
13'b1100011010110: edge_mask_reg_512p3[228] <= 1'b1;
 		default: edge_mask_reg_512p3[228] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[229] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[230] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[231] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[232] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101111001,
13'b100011001000,
13'b100011001001,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b110011011000,
13'b110011011001,
13'b110011101000,
13'b110011101001,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101001000,
13'b110101001001,
13'b110101011000,
13'b110101011001,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1011011110100,
13'b1011011110101,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011101000011,
13'b1100100000100,
13'b1100100000101,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100010101,
13'b1100100010110,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100100110101,
13'b1100101000011,
13'b1101100010010,
13'b1101100010011,
13'b1101100010100,
13'b1101100100010,
13'b1101100100011,
13'b1101100100100,
13'b1101100100101,
13'b1101100100110,
13'b1101100110011,
13'b1101100110100: edge_mask_reg_512p3[233] <= 1'b1;
 		default: edge_mask_reg_512p3[233] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b101011011000,
13'b101011011001,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b110011101000,
13'b110011101001,
13'b110011111000,
13'b110011111001,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110011000,
13'b110110011001,
13'b111011110110,
13'b111011110111,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000101,
13'b111110000110,
13'b1000011110110,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000100,
13'b1001110000101,
13'b1010100000100,
13'b1010100000101,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000010,
13'b1010110000100,
13'b1010110000101,
13'b1011100000100,
13'b1011100000101,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1100100000101,
13'b1100100010011,
13'b1100100010100,
13'b1100100010101,
13'b1100100010110,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100100110101,
13'b1100100110110,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101010101,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110010,
13'b1100101110100,
13'b1100101110101,
13'b1101100100010,
13'b1101100100011,
13'b1101100100100,
13'b1101100100101,
13'b1101100100110,
13'b1101100110010,
13'b1101100110011,
13'b1101100110100,
13'b1101100110101,
13'b1101101000010,
13'b1101101000011,
13'b1101101010011: edge_mask_reg_512p3[234] <= 1'b1;
 		default: edge_mask_reg_512p3[234] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001001,
13'b101111001010,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100101,
13'b110110100110,
13'b111011110111,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b1000011110110,
13'b1000011110111,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1010011110101,
13'b1010011110110,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010100,
13'b1010110010101,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110010,
13'b1011101110100,
13'b1011101110101,
13'b1100100000011,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100010011,
13'b1100100010100,
13'b1100100010101,
13'b1100100010110,
13'b1100100100011,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100110011,
13'b1100100110100,
13'b1100100110101,
13'b1100100110110,
13'b1100101000011: edge_mask_reg_512p3[235] <= 1'b1;
 		default: edge_mask_reg_512p3[235] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100101,
13'b101100110,
13'b101100111,
13'b1101110101,
13'b1101110110,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b101110000101,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111100000,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111110000,
13'b1010111110001,
13'b1010111110010,
13'b1010111110011,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111010000,
13'b1011111010001,
13'b1011111010010,
13'b1011111100000,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111110000,
13'b1011111110001,
13'b1011111110010,
13'b1011111110011,
13'b1100111000000,
13'b1100111000001,
13'b1100111010000,
13'b1100111010001,
13'b1100111010010,
13'b1100111100000,
13'b1100111100001,
13'b1100111100010,
13'b1100111110000,
13'b1100111110001,
13'b1100111110010,
13'b1100111110011,
13'b1101111100001,
13'b1101111100010,
13'b1101111110000,
13'b1101111110001,
13'b1101111110010: edge_mask_reg_512p3[236] <= 1'b1;
 		default: edge_mask_reg_512p3[236] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11011101,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11101101,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b11111101,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100001101,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100011101,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100101101,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011011101,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011101101,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1011111101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100001101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100011101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100101101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111010,
13'b1101111011,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101000110,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111010,
13'b10101111011,
13'b11001101010,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101000110,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101010,
13'b11101101011,
13'b100001111001,
13'b100001111010,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111010,
13'b100100111011,
13'b101010001010,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010011010,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111010,
13'b101010111011,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001010,
13'b101011001011,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011010,
13'b101011011011,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101010,
13'b101011101011,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111010,
13'b101011111011,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110101,
13'b101100110110,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100010011,
13'b110100010100,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111100000011,
13'b111100000100,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110011,
13'b1001011000011,
13'b1001011010011: edge_mask_reg_512p3[237] <= 1'b1;
 		default: edge_mask_reg_512p3[237] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101000111,
13'b110101001000,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101100101,
13'b111101100110,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1001101100100,
13'b1001101100101,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1011101100011,
13'b1011101100100,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1100101100011,
13'b1100101110001,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100110000001,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111010011,
13'b1100111010100,
13'b1101101110001,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1101110000001,
13'b1101110000010,
13'b1101110000011,
13'b1101110000100,
13'b1101110010001,
13'b1101110010010,
13'b1101110010011,
13'b1101110010100,
13'b1101110100001,
13'b1101110100010,
13'b1101110100011,
13'b1101110100100,
13'b1101110110001,
13'b1101110110010,
13'b1101110110011,
13'b1101110110100,
13'b1101111000001,
13'b1101111000010,
13'b1101111000011,
13'b1110101110001,
13'b1110101110010,
13'b1110110000001,
13'b1110110000010,
13'b1110110010001,
13'b1110110010010,
13'b1110110010011,
13'b1110110100001,
13'b1110110100010,
13'b1110110100011,
13'b1110110110001,
13'b1110110110010,
13'b1110110110011,
13'b1110111000001,
13'b1110111000010,
13'b1110111000011: edge_mask_reg_512p3[238] <= 1'b1;
 		default: edge_mask_reg_512p3[238] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110000110,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b1000110000101,
13'b1000110000110,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111010011,
13'b1100111010100,
13'b1101110010010,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1101110100001,
13'b1101110100010,
13'b1101110100011,
13'b1101110100100,
13'b1101110100101,
13'b1101110110001,
13'b1101110110010,
13'b1101110110011,
13'b1101110110100,
13'b1101111000001,
13'b1101111000010,
13'b1101111000011,
13'b1110110010010,
13'b1110110100010,
13'b1110110100011,
13'b1110110110001,
13'b1110110110010,
13'b1110110110011,
13'b1110111000001,
13'b1110111000010,
13'b1110111000011: edge_mask_reg_512p3[239] <= 1'b1;
 		default: edge_mask_reg_512p3[239] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101110111,
13'b101101111000,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001110010101,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111110001,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111010000,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100000,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111110000,
13'b1011111110001,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111010000,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111100000,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111110000,
13'b1100111110001,
13'b1100111110010,
13'b1100111110011,
13'b1100111110100,
13'b1101110100001,
13'b1101110100010,
13'b1101110100011,
13'b1101110100100,
13'b1101110110001,
13'b1101110110010,
13'b1101110110011,
13'b1101110110100,
13'b1101111000001,
13'b1101111000010,
13'b1101111000011,
13'b1101111000100,
13'b1101111010000,
13'b1101111010001,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1101111100000,
13'b1101111100001,
13'b1101111100010,
13'b1101111100011,
13'b1101111110000,
13'b1101111110001,
13'b1101111110010,
13'b1101111110011,
13'b1110110100001,
13'b1110110100010,
13'b1110110110001,
13'b1110110110010,
13'b1110111000001,
13'b1110111000010,
13'b1110111000011,
13'b1110111010001,
13'b1110111010010,
13'b1110111100000,
13'b1110111100001,
13'b1110111100010,
13'b1110111110000,
13'b1110111110001: edge_mask_reg_512p3[240] <= 1'b1;
 		default: edge_mask_reg_512p3[240] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[241] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100111,
13'b11100101000,
13'b100000110111,
13'b100000111000,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010010,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100001,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100111,
13'b100100101000,
13'b101000110111,
13'b101000111000,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100111,
13'b101100101000,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010111,
13'b110100011000,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110111,
13'b111001111000,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000111,
13'b111010001000,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010111,
13'b111010011000,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100111,
13'b111010101000,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000000,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b1000001110000,
13'b1000001110010,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010010000,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010100000,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010110000,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000000,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010000,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1001010000000,
13'b1001010010000,
13'b1001010010001,
13'b1001010100000,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010110000,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1010010100000,
13'b1010010100001,
13'b1010010110000,
13'b1010010110001,
13'b1010011000000,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011110010,
13'b1010011110011,
13'b1011010110000,
13'b1011010110001,
13'b1011011000000,
13'b1011011000001,
13'b1011011010000,
13'b1011011010001,
13'b1011011100000,
13'b1011011100001,
13'b1100011010000,
13'b1100011010001,
13'b1100011100000: edge_mask_reg_512p3[242] <= 1'b1;
 		default: edge_mask_reg_512p3[242] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b100011111000,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110111,
13'b100110111000,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100111,
13'b110110101000,
13'b111100100111,
13'b111100101000,
13'b111100110111,
13'b111100111000,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110110,
13'b1000101110111,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1010100100111,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1011100100110,
13'b1011100100111,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110101,
13'b1011101110110,
13'b1011101110111,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100101,
13'b1100101100110,
13'b1100101100111,
13'b1100101110101,
13'b1100101110110,
13'b1100101110111,
13'b1101100100111,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101010100,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101100100,
13'b1101101100101,
13'b1101101100110,
13'b1101101100111,
13'b1101101110101,
13'b1101101110110,
13'b1101101110111,
13'b1110100110101,
13'b1110100110110,
13'b1110100110111,
13'b1110101000101,
13'b1110101000110,
13'b1110101000111,
13'b1110101010100,
13'b1110101010101,
13'b1110101010110,
13'b1110101010111,
13'b1110101100100,
13'b1110101100101,
13'b1110101100110,
13'b1110101100111,
13'b1110101110101,
13'b1110101110110,
13'b1111100110101,
13'b1111100110110,
13'b1111100110111,
13'b1111101000101,
13'b1111101000110,
13'b1111101000111,
13'b1111101010100,
13'b1111101010101,
13'b1111101010110,
13'b1111101010111,
13'b1111101100011,
13'b1111101100100,
13'b1111101100101,
13'b1111101100110,
13'b1111101100111,
13'b1111101110101,
13'b1111101110110: edge_mask_reg_512p3[243] <= 1'b1;
 		default: edge_mask_reg_512p3[243] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111101010110,
13'b111101010111,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100111,
13'b111111101000,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000110,
13'b1000110000111,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010111,
13'b1001111011000,
13'b1001111100111,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110110,
13'b1010110110111,
13'b1010110111000,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111010111,
13'b1010111011000,
13'b1010111100111,
13'b1011101010101,
13'b1011101010110,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1011101110101,
13'b1011101110110,
13'b1011101110111,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110110110,
13'b1011110110111,
13'b1011110111000,
13'b1011111000110,
13'b1011111000111,
13'b1011111001000,
13'b1011111010111,
13'b1011111011000,
13'b1011111100111,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1100101100100,
13'b1100101100101,
13'b1100101100110,
13'b1100101100111,
13'b1100101110100,
13'b1100101110101,
13'b1100101110110,
13'b1100101110111,
13'b1100110000101,
13'b1100110000110,
13'b1100110000111,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1100110100110,
13'b1100110100111,
13'b1100110101000,
13'b1100110110110,
13'b1100110110111,
13'b1100110111000,
13'b1100111000110,
13'b1100111000111,
13'b1100111001000,
13'b1100111010111,
13'b1100111011000,
13'b1101101010100,
13'b1101101010101,
13'b1101101010110,
13'b1101101100011,
13'b1101101100100,
13'b1101101100101,
13'b1101101100110,
13'b1101101110011,
13'b1101101110100,
13'b1101101110101,
13'b1101101110110,
13'b1101101110111,
13'b1101110000100,
13'b1101110000101,
13'b1101110000110,
13'b1101110000111,
13'b1101110010101,
13'b1101110010110,
13'b1101110010111,
13'b1101110100101,
13'b1101110100110,
13'b1101110100111,
13'b1101110101000,
13'b1101110110110,
13'b1101110110111,
13'b1101110111000,
13'b1101111000110,
13'b1101111000111,
13'b1101111001000,
13'b1101111010111,
13'b1101111011000,
13'b1110101010100,
13'b1110101010101,
13'b1110101010110,
13'b1110101100011,
13'b1110101100100,
13'b1110101100101,
13'b1110101100110,
13'b1110101110011,
13'b1110101110100,
13'b1110101110101,
13'b1110101110110,
13'b1110101110111,
13'b1110110000011,
13'b1110110000100,
13'b1110110000101,
13'b1110110000110,
13'b1110110000111,
13'b1110110010100,
13'b1110110010101,
13'b1110110010110,
13'b1110110010111,
13'b1110110100100,
13'b1110110100101,
13'b1110110100110,
13'b1110110100111,
13'b1110110101000,
13'b1110110110101,
13'b1110110110110,
13'b1110110110111,
13'b1110110111000,
13'b1110111000110,
13'b1110111000111,
13'b1110111001000,
13'b1110111010110,
13'b1110111010111,
13'b1110111011000,
13'b1111101010101,
13'b1111101010110,
13'b1111101100011,
13'b1111101100100,
13'b1111101100101,
13'b1111101100110,
13'b1111101110011,
13'b1111101110100,
13'b1111101110101,
13'b1111101110110,
13'b1111101110111,
13'b1111110000011,
13'b1111110000100,
13'b1111110000101,
13'b1111110000110,
13'b1111110000111,
13'b1111110010011,
13'b1111110010100,
13'b1111110010101,
13'b1111110010110,
13'b1111110010111,
13'b1111110100100,
13'b1111110100101,
13'b1111110100110,
13'b1111110100111,
13'b1111110101000,
13'b1111110110100,
13'b1111110110101,
13'b1111110110110,
13'b1111110110111,
13'b1111110111000,
13'b1111111000101,
13'b1111111000110,
13'b1111111000111,
13'b1111111001000,
13'b1111111010110,
13'b1111111010111,
13'b1111111011000: edge_mask_reg_512p3[244] <= 1'b1;
 		default: edge_mask_reg_512p3[244] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10101000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b100000110000,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000000,
13'b100001000001,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010000,
13'b100001010010,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100000,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110011,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1011000100010,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001010000,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001100000,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1100001000010,
13'b1100001000011,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1100001100010,
13'b1100001100011: edge_mask_reg_512p3[245] <= 1'b1;
 		default: edge_mask_reg_512p3[245] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100011111000,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110011000,
13'b110110011001,
13'b110110101001,
13'b111100100111,
13'b111100101000,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101110111,
13'b1000101111000,
13'b1000101111001,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110111,
13'b1001101111000,
13'b1001101111001,
13'b1001110000111,
13'b1001110001000,
13'b1001110001001,
13'b1010100100111,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010101111001,
13'b1010110000111,
13'b1010110001000,
13'b1010110001001,
13'b1011100100110,
13'b1011100100111,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1011110000111,
13'b1011110001000,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1101100100111,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1110100110101,
13'b1110100110110,
13'b1110100110111,
13'b1110101000101,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101010101,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110110000111,
13'b1110110001000,
13'b1111100110101,
13'b1111100110110,
13'b1111100110111,
13'b1111101000101,
13'b1111101000110,
13'b1111101000111,
13'b1111101010101,
13'b1111101010110,
13'b1111101010111,
13'b1111101011000,
13'b1111101100110,
13'b1111101100111,
13'b1111101101000,
13'b1111101110110,
13'b1111101110111,
13'b1111101111000: edge_mask_reg_512p3[246] <= 1'b1;
 		default: edge_mask_reg_512p3[246] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101000,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b110100101000,
13'b110100101001,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110001000,
13'b110110001001,
13'b110110011000,
13'b110110011001,
13'b110110101001,
13'b111100111000,
13'b111100111001,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101110111,
13'b1000101111000,
13'b1000101111001,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1001100111000,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110111,
13'b1001101111000,
13'b1001101111001,
13'b1001110000111,
13'b1001110001000,
13'b1001110001001,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101010111,
13'b1010101011000,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110111,
13'b1010101111000,
13'b1010101111001,
13'b1010110000111,
13'b1010110001000,
13'b1010110001001,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110111,
13'b1011101111000,
13'b1011110000111,
13'b1011110001000,
13'b1100100110111,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100110000111,
13'b1100110001000,
13'b1101100110111,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101110000111,
13'b1101110001000,
13'b1110100110111,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110110000111,
13'b1110110001000,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111,
13'b1111101011000,
13'b1111101100110,
13'b1111101100111,
13'b1111101101000,
13'b1111101110110,
13'b1111101110111,
13'b1111101111000: edge_mask_reg_512p3[247] <= 1'b1;
 		default: edge_mask_reg_512p3[247] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110100101,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001110100101,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010110100100,
13'b1010110100101,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111100110,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110,
13'b1101110110011,
13'b1101110110100,
13'b1101111000010,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1101111010101,
13'b1101111100010,
13'b1101111100011,
13'b1101111100100,
13'b1101111100101,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1101111110110,
13'b1110110110010,
13'b1110110110011,
13'b1110111000010,
13'b1110111000011,
13'b1110111000100,
13'b1110111010010,
13'b1110111010011,
13'b1110111010100,
13'b1110111100010,
13'b1110111100011,
13'b1110111100100,
13'b1110111100101,
13'b1110111110010,
13'b1110111110011,
13'b1110111110100,
13'b1110111110101,
13'b1111110110010,
13'b1111110110011,
13'b1111111000010,
13'b1111111000011,
13'b1111111000100,
13'b1111111010010,
13'b1111111010011,
13'b1111111010100,
13'b1111111100010,
13'b1111111100011,
13'b1111111100100,
13'b1111111110010,
13'b1111111110011,
13'b1111111110100,
13'b1111111110101: edge_mask_reg_512p3[248] <= 1'b1;
 		default: edge_mask_reg_512p3[248] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[249] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[250] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101110111,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101110111,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111100000,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111110000,
13'b1010111110001,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1011110100010,
13'b1011110100011,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111010000,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111100000,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111110001,
13'b1011111110010,
13'b1011111110011,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111010000,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111100010,
13'b1100111100011: edge_mask_reg_512p3[251] <= 1'b1;
 		default: edge_mask_reg_512p3[251] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101100111,
13'b100101101000,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101100111,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110000,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110000011,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1010110010010,
13'b1010110010011,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111100000,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111110000,
13'b1010111110001,
13'b1010111110010,
13'b1010111110011,
13'b1011110010010,
13'b1011110010011,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111010010,
13'b1011111010011,
13'b1011111100010,
13'b1011111100011,
13'b1011111110010,
13'b1011111110011: edge_mask_reg_512p3[252] <= 1'b1;
 		default: edge_mask_reg_512p3[252] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101110111,
13'b100101111000,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101110111,
13'b101101111000,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010000,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110000111,
13'b110110001000,
13'b110110010010,
13'b110110010011,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110010010,
13'b111110010011,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110111,
13'b111110111000,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100111,
13'b111111101000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1001110110010,
13'b1001110110011,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011: edge_mask_reg_512p3[253] <= 1'b1;
 		default: edge_mask_reg_512p3[253] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100110,
13'b101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100110000110,
13'b100110000111,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101110000110,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100001,
13'b101110100010,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111110100000,
13'b111110100001,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000110,
13'b111111000111,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010110,
13'b111111010111,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100110,
13'b111111100111,
13'b1000110110000,
13'b1000110110001,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1001111010001,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010: edge_mask_reg_512p3[254] <= 1'b1;
 		default: edge_mask_reg_512p3[254] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010111,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000000,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010000,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100000,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110000,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100100110101,
13'b100100110110,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101100110101,
13'b101100110110,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111101100000,
13'b111101110000,
13'b111101110001,
13'b111101110101,
13'b111101110110,
13'b111110000000,
13'b111110000001,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110110,
13'b111110110111,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000110,
13'b111111000111,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b1000110100000,
13'b1000110100001,
13'b1000110110000,
13'b1000110110001,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111010000,
13'b1000111010001: edge_mask_reg_512p3[255] <= 1'b1;
 		default: edge_mask_reg_512p3[255] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000000,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110000,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000101,
13'b101111000110,
13'b110011100110,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000001,
13'b110100000010,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110111000101,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010110,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100110,
13'b111100100111,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110110,
13'b111100110111,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110101,
13'b111101110110,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000101,
13'b111110000110,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010101,
13'b111110010110,
13'b111110100000,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000110000000,
13'b1000110000001,
13'b1000110010000,
13'b1001100000000,
13'b1001100000001,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100100000,
13'b1001100100001,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101010000,
13'b1001101010001,
13'b1001101100000,
13'b1001101100001,
13'b1010100010000,
13'b1010100010001,
13'b1010100100000,
13'b1010100100001,
13'b1010100110000,
13'b1010100110001,
13'b1010101000000,
13'b1010101000001: edge_mask_reg_512p3[256] <= 1'b1;
 		default: edge_mask_reg_512p3[256] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10010110111,
13'b10010111000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110111000,
13'b11110111001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110111000,
13'b100110111001,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110111000,
13'b101110111001,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b111011100110,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000101,
13'b111110000110,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1010011100011,
13'b1010011100100,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1100011110001,
13'b1100011110010,
13'b1100011110011,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100000100,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100110000100,
13'b1101011110001,
13'b1101011110010,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100100001,
13'b1101100100010,
13'b1101100100011,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101010100,
13'b1101101100010,
13'b1101101100011,
13'b1101101100100,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1110100000010,
13'b1110100010010,
13'b1110100010011,
13'b1110100100010,
13'b1110100100011,
13'b1110100110010,
13'b1110100110011,
13'b1110101000010,
13'b1110101000011,
13'b1110101010010,
13'b1110101010011,
13'b1110101100010,
13'b1110101100011,
13'b1110101110010,
13'b1110101110011: edge_mask_reg_512p3[257] <= 1'b1;
 		default: edge_mask_reg_512p3[257] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100000111,
13'b1100001000,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011000,
13'b100100011001,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000101,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101000101,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1011101000011,
13'b1011101000100,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1101101010010,
13'b1101101010011,
13'b1101101100010,
13'b1101101100011,
13'b1101101100100,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1101110000010,
13'b1101110000011,
13'b1101110000100,
13'b1101110010010,
13'b1101110010011,
13'b1101110010100,
13'b1101110100010,
13'b1101110100011,
13'b1101110100100,
13'b1101110110010,
13'b1101110110011,
13'b1101110110100,
13'b1101111000010,
13'b1101111000011,
13'b1101111000100,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1110101010010,
13'b1110101010011,
13'b1110101100010,
13'b1110101100011,
13'b1110101110010,
13'b1110101110011,
13'b1110110000010,
13'b1110110000011,
13'b1110110010010,
13'b1110110010011,
13'b1110110010100,
13'b1110110100010,
13'b1110110100011,
13'b1110110100100,
13'b1110110110010,
13'b1110110110011,
13'b1110110110100,
13'b1110111000010,
13'b1110111000011,
13'b1110111000100,
13'b1110111010010,
13'b1110111010011,
13'b1110111010100,
13'b1111101110011,
13'b1111110000010,
13'b1111110000011,
13'b1111110010010,
13'b1111110010011,
13'b1111110100010,
13'b1111110100011,
13'b1111110110010,
13'b1111110110011,
13'b1111111000010,
13'b1111111000011,
13'b1111111000100,
13'b1111111010010,
13'b1111111010011: edge_mask_reg_512p3[258] <= 1'b1;
 		default: edge_mask_reg_512p3[258] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b100100011000,
13'b100100011001,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000101,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011101110111,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101100110,
13'b1100101100111,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100101110110,
13'b1100101110111,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110000111,
13'b1101101000101,
13'b1101101000110,
13'b1101101010010,
13'b1101101010011,
13'b1101101010100,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101100010,
13'b1101101100011,
13'b1101101100100,
13'b1101101100101,
13'b1101101100110,
13'b1101101100111,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1101101110101,
13'b1101101110110,
13'b1101101110111,
13'b1101110000101,
13'b1101110000110,
13'b1110101010010,
13'b1110101010011,
13'b1110101010100,
13'b1110101010101,
13'b1110101010110,
13'b1110101100010,
13'b1110101100011,
13'b1110101100100,
13'b1110101100101,
13'b1110101100110,
13'b1110101110010,
13'b1110101110011,
13'b1110101110100,
13'b1110101110101,
13'b1110101110110,
13'b1111101010011,
13'b1111101010100,
13'b1111101010101,
13'b1111101010110,
13'b1111101100011,
13'b1111101100100,
13'b1111101100101,
13'b1111101100110,
13'b1111101110011,
13'b1111101110100,
13'b1111101110101,
13'b1111101110110: edge_mask_reg_512p3[259] <= 1'b1;
 		default: edge_mask_reg_512p3[259] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1100000111,
13'b1100001000,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100100011000,
13'b100100011001,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000101,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101000101,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010111,
13'b111111011000,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010110111000,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111010110,
13'b1010111010111,
13'b1010111011000,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010101,
13'b1011111010110,
13'b1011111010111,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101010101,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100101110110,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1100110100100,
13'b1100110100101,
13'b1100110100110,
13'b1100110100111,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111010101,
13'b1100111010110,
13'b1100111010111,
13'b1101101010010,
13'b1101101010011,
13'b1101101100010,
13'b1101101100011,
13'b1101101100100,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1101101110101,
13'b1101110000010,
13'b1101110000011,
13'b1101110000100,
13'b1101110000101,
13'b1101110000110,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1101110010110,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1101110100111,
13'b1101110110100,
13'b1101110110101,
13'b1101110110110,
13'b1101110110111,
13'b1101111000101,
13'b1101111000110,
13'b1101111000111,
13'b1101111010110,
13'b1110101010010,
13'b1110101010011,
13'b1110101100010,
13'b1110101100011,
13'b1110101100100,
13'b1110101110010,
13'b1110101110011,
13'b1110101110100,
13'b1110101110101,
13'b1110110000010,
13'b1110110000011,
13'b1110110000100,
13'b1110110000101,
13'b1110110010011,
13'b1110110010100,
13'b1110110010101,
13'b1110110010110,
13'b1110110100011,
13'b1110110100100,
13'b1110110100101,
13'b1110110100110,
13'b1110110110100,
13'b1110110110101,
13'b1110110110110,
13'b1110110110111,
13'b1110111000101,
13'b1110111000110,
13'b1111101100011,
13'b1111101110011,
13'b1111101110100,
13'b1111110000011,
13'b1111110000100,
13'b1111110000101,
13'b1111110010011,
13'b1111110010100,
13'b1111110010101,
13'b1111110010110,
13'b1111110100100,
13'b1111110100101,
13'b1111110100110,
13'b1111110110100,
13'b1111110110101,
13'b1111110110110,
13'b1111111000101,
13'b1111111000110: edge_mask_reg_512p3[260] <= 1'b1;
 		default: edge_mask_reg_512p3[260] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110111000,
13'b11110111001,
13'b100011000111,
13'b100011001000,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110111000,
13'b100110111001,
13'b101011000111,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110111000,
13'b101110111001,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000101,
13'b111110000110,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1100011110010,
13'b1100011110011,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100110000100,
13'b1101100000000,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100100001,
13'b1101100100010,
13'b1101100100011,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101010100,
13'b1101101100010,
13'b1101101100011,
13'b1101101100100,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1110100000001,
13'b1110100000010,
13'b1110100010001,
13'b1110100010010,
13'b1110100100001,
13'b1110100100010,
13'b1110100100011,
13'b1110100110001,
13'b1110100110010,
13'b1110100110011,
13'b1110101000001,
13'b1110101000010,
13'b1110101000011,
13'b1110101010010,
13'b1110101010011,
13'b1110101100010,
13'b1110101100011,
13'b1110101110010,
13'b1110101110011,
13'b1111100010001,
13'b1111100010010,
13'b1111100100010,
13'b1111100110010,
13'b1111101000010,
13'b1111101010010: edge_mask_reg_512p3[261] <= 1'b1;
 		default: edge_mask_reg_512p3[261] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110101,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011000110,
13'b10011000111,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b101011010110,
13'b101011010111,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100101,
13'b101110100110,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100101,
13'b110110100110,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1001011110100,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1101100000001,
13'b1101100000010,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100100000,
13'b1101100100001,
13'b1101100100010,
13'b1101100100011,
13'b1101100100100,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101100110100,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101000100,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101010100,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1101101100100,
13'b1101101110001,
13'b1101101110010,
13'b1101101110011,
13'b1110100000000,
13'b1110100000001,
13'b1110100010000,
13'b1110100010001,
13'b1110100010010,
13'b1110100100000,
13'b1110100100001,
13'b1110100100010,
13'b1110100110000,
13'b1110100110001,
13'b1110100110010,
13'b1110100110011,
13'b1110101000000,
13'b1110101000001,
13'b1110101000010,
13'b1110101000011,
13'b1110101000100,
13'b1110101010000,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101010100,
13'b1110101100000,
13'b1110101100001,
13'b1110101100010,
13'b1110101100011,
13'b1110101100100,
13'b1110101110001,
13'b1110101110010,
13'b1110101110011,
13'b1111100010001,
13'b1111100010010,
13'b1111100100000,
13'b1111100100001,
13'b1111100100010,
13'b1111100110000,
13'b1111100110001,
13'b1111100110010,
13'b1111101000000,
13'b1111101000001,
13'b1111101000010,
13'b1111101010000,
13'b1111101010001,
13'b1111101010010,
13'b1111101100000,
13'b1111101100001,
13'b1111101100010,
13'b1111101110001,
13'b1111101110010: edge_mask_reg_512p3[262] <= 1'b1;
 		default: edge_mask_reg_512p3[262] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100110,
13'b100100111,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100110110,
13'b1100110111,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101000110,
13'b100101000111,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101000110,
13'b101101000111,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101010110,
13'b110101010111,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100110000001,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111010110,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111100110,
13'b1100111110010,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110,
13'b1101101110011,
13'b1101101110100,
13'b1101110000001,
13'b1101110000010,
13'b1101110000011,
13'b1101110000100,
13'b1101110010001,
13'b1101110010010,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1101110100001,
13'b1101110100010,
13'b1101110100011,
13'b1101110100100,
13'b1101110100101,
13'b1101110110001,
13'b1101110110010,
13'b1101110110011,
13'b1101110110100,
13'b1101110110101,
13'b1101111000001,
13'b1101111000010,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111010001,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1101111010101,
13'b1101111100010,
13'b1101111100011,
13'b1101111100100,
13'b1101111100101,
13'b1101111110010,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1110101110011,
13'b1110101110100,
13'b1110110000001,
13'b1110110000010,
13'b1110110000011,
13'b1110110000100,
13'b1110110010001,
13'b1110110010010,
13'b1110110010011,
13'b1110110010100,
13'b1110110100001,
13'b1110110100010,
13'b1110110100011,
13'b1110110100100,
13'b1110110100101,
13'b1110110110001,
13'b1110110110010,
13'b1110110110011,
13'b1110110110100,
13'b1110110110101,
13'b1110111000001,
13'b1110111000010,
13'b1110111000011,
13'b1110111000100,
13'b1110111000101,
13'b1110111010010,
13'b1110111010011,
13'b1110111010100,
13'b1110111010101,
13'b1110111100010,
13'b1110111100011,
13'b1110111100100,
13'b1110111100101,
13'b1110111110010,
13'b1110111110011,
13'b1110111110100,
13'b1110111110101,
13'b1111110010001,
13'b1111110010010,
13'b1111110100001,
13'b1111110100010,
13'b1111110110001,
13'b1111110110010,
13'b1111111000010,
13'b1111111000011,
13'b1111111010010,
13'b1111111010011,
13'b1111111100010,
13'b1111111100011,
13'b1111111110010,
13'b1111111110011: edge_mask_reg_512p3[263] <= 1'b1;
 		default: edge_mask_reg_512p3[263] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100110,
13'b101100111,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101110110,
13'b100101110111,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101110110,
13'b101101110111,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110000110,
13'b110110000111,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100000,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111010000,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100000,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010000,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111100000,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111110001,
13'b1100111110010,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110,
13'b1101111000010,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111010000,
13'b1101111010001,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1101111010101,
13'b1101111100000,
13'b1101111100001,
13'b1101111100010,
13'b1101111100011,
13'b1101111100100,
13'b1101111100101,
13'b1101111110001,
13'b1101111110010,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1110111010100,
13'b1110111010101,
13'b1110111100001,
13'b1110111100010,
13'b1110111100011,
13'b1110111100100,
13'b1110111100101,
13'b1110111110001,
13'b1110111110010,
13'b1110111110011,
13'b1110111110100,
13'b1110111110101,
13'b1111111110010,
13'b1111111110011: edge_mask_reg_512p3[264] <= 1'b1;
 		default: edge_mask_reg_512p3[264] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000110,
13'b101000111,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101010110,
13'b1101010111,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101100110,
13'b101101100111,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110000011,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110000010,
13'b1000110000011,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010000,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001110000001,
13'b1001110000010,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100000,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111010000,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100000,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010000,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111100000,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111110001,
13'b1100111110010,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111010000,
13'b1101111010001,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1101111010101,
13'b1101111100001,
13'b1101111100010,
13'b1101111100011,
13'b1101111100100,
13'b1101111100101,
13'b1101111110001,
13'b1101111110010,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1110111010100,
13'b1110111010101,
13'b1110111100001,
13'b1110111100010,
13'b1110111100011,
13'b1110111100100,
13'b1110111100101,
13'b1110111110001,
13'b1110111110010,
13'b1110111110011,
13'b1110111110100,
13'b1110111110101,
13'b1111111110010,
13'b1111111110011: edge_mask_reg_512p3[265] <= 1'b1;
 		default: edge_mask_reg_512p3[265] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100011000,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100111000,
13'b100100111001,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100111000,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101011000,
13'b110101011001,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1100101100100,
13'b1100101100101,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110010110,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110100110,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100110110110,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111000110,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111010110,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111100110,
13'b1100111110010,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1101101110101,
13'b1101110000010,
13'b1101110000011,
13'b1101110000100,
13'b1101110000101,
13'b1101110010010,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1101110100010,
13'b1101110100011,
13'b1101110100100,
13'b1101110100101,
13'b1101110110010,
13'b1101110110011,
13'b1101110110100,
13'b1101110110101,
13'b1101111000010,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1101111010101,
13'b1101111100010,
13'b1101111100011,
13'b1101111100100,
13'b1101111100101,
13'b1101111110010,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1110110000010,
13'b1110110000011,
13'b1110110010010,
13'b1110110010011,
13'b1110110100010,
13'b1110110100011,
13'b1110110110010,
13'b1110110110011,
13'b1110111000010,
13'b1110111000011,
13'b1110111000100,
13'b1110111000101,
13'b1110111010010,
13'b1110111010011,
13'b1110111010100,
13'b1110111010101,
13'b1110111100010,
13'b1110111100011,
13'b1110111100100,
13'b1110111100101,
13'b1110111110010,
13'b1110111110011,
13'b1110111110100,
13'b1110111110101,
13'b1111111000010,
13'b1111111010010,
13'b1111111010011,
13'b1111111100010,
13'b1111111100011,
13'b1111111110010,
13'b1111111110011: edge_mask_reg_512p3[266] <= 1'b1;
 		default: edge_mask_reg_512p3[266] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100110110,
13'b100110111,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101000110,
13'b1101000111,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101101010110,
13'b101101010111,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1100110000010,
13'b1100110000011,
13'b1100110010000,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110100000,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1100110110000,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111100110,
13'b1100111110001,
13'b1100111110010,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110,
13'b1101110010010,
13'b1101110010011,
13'b1101110100000,
13'b1101110100001,
13'b1101110100010,
13'b1101110100011,
13'b1101110100100,
13'b1101110110000,
13'b1101110110001,
13'b1101110110010,
13'b1101110110011,
13'b1101110110100,
13'b1101111000000,
13'b1101111000001,
13'b1101111000010,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111010001,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1101111010101,
13'b1101111100001,
13'b1101111100010,
13'b1101111100011,
13'b1101111100100,
13'b1101111100101,
13'b1101111110001,
13'b1101111110010,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1110111000001,
13'b1110111000010,
13'b1110111010001,
13'b1110111010010,
13'b1110111010011,
13'b1110111010100,
13'b1110111010101,
13'b1110111100001,
13'b1110111100010,
13'b1110111100011,
13'b1110111100100,
13'b1110111100101,
13'b1110111110010,
13'b1110111110011,
13'b1110111110100,
13'b1110111110101,
13'b1111111100010,
13'b1111111110010,
13'b1111111110011: edge_mask_reg_512p3[267] <= 1'b1;
 		default: edge_mask_reg_512p3[267] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001111000110,
13'b1001111000111,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010111000110,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1011111000101,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1011111110111,
13'b1100111000101,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111010110,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111100110,
13'b1100111110010,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110,
13'b1101111010011,
13'b1101111010100,
13'b1101111010101,
13'b1101111010110,
13'b1101111100010,
13'b1101111100011,
13'b1101111100100,
13'b1101111100101,
13'b1101111100110,
13'b1101111110010,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1101111110110,
13'b1110111010100,
13'b1110111010101,
13'b1110111100010,
13'b1110111100011,
13'b1110111100100,
13'b1110111100101,
13'b1110111110010,
13'b1110111110011,
13'b1110111110100,
13'b1110111110101,
13'b1110111110110,
13'b1111111100010,
13'b1111111100011,
13'b1111111110010,
13'b1111111110011,
13'b1111111110100: edge_mask_reg_512p3[268] <= 1'b1;
 		default: edge_mask_reg_512p3[268] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100111,
13'b11011101000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100111,
13'b100011101000,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100111,
13'b101011101000,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010111,
13'b110011011000,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110111,
13'b111010111000,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010001001,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010111000,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010001001,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010111000,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001010101,
13'b1010001010110,
13'b1010001010111,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001101000,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010001001,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010111000,
13'b1011000010100,
13'b1011000010101,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001000111,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001010111,
13'b1011001100101,
13'b1011001100110,
13'b1011001100111,
13'b1011001101000,
13'b1011001110110,
13'b1011001110111,
13'b1011001111000,
13'b1011010000110,
13'b1011010000111,
13'b1011010001000,
13'b1011010001001,
13'b1011010010111,
13'b1011010011000,
13'b1011010011001,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010111000,
13'b1011010111001,
13'b1100000010011,
13'b1100000010100,
13'b1100000010101,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000100110,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100000110110,
13'b1100001000100,
13'b1100001000101,
13'b1100001000110,
13'b1100001000111,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001010111,
13'b1100001100101,
13'b1100001100110,
13'b1100001100111,
13'b1100001101000,
13'b1100001110110,
13'b1100001110111,
13'b1100001111000,
13'b1100010000110,
13'b1100010000111,
13'b1100010001000,
13'b1100010001001,
13'b1100010010111,
13'b1100010011000,
13'b1100010011001,
13'b1100010100111,
13'b1100010101000,
13'b1100010101001,
13'b1100010111000,
13'b1100010111001,
13'b1101000010011,
13'b1101000010100,
13'b1101000010101,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000100110,
13'b1101000110010,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101000110110,
13'b1101001000010,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001000110,
13'b1101001000111,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001010110,
13'b1101001010111,
13'b1101001100101,
13'b1101001100110,
13'b1101001100111,
13'b1101001101000,
13'b1101001110101,
13'b1101001110110,
13'b1101001110111,
13'b1101001111000,
13'b1101001111001,
13'b1101010000110,
13'b1101010000111,
13'b1101010001000,
13'b1101010001001,
13'b1101010010111,
13'b1101010011000,
13'b1101010011001,
13'b1101010011010,
13'b1101010100111,
13'b1101010101000,
13'b1101010101001,
13'b1101010101010,
13'b1101010111000,
13'b1101010111001,
13'b1110000010011,
13'b1110000010100,
13'b1110000010101,
13'b1110000100010,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000110010,
13'b1110000110011,
13'b1110000110100,
13'b1110000110101,
13'b1110000110110,
13'b1110001000010,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1110001000110,
13'b1110001000111,
13'b1110001010010,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001010110,
13'b1110001010111,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001100110,
13'b1110001100111,
13'b1110001101000,
13'b1110001110100,
13'b1110001110101,
13'b1110001110110,
13'b1110001110111,
13'b1110001111000,
13'b1110001111001,
13'b1110010000101,
13'b1110010000110,
13'b1110010000111,
13'b1110010001000,
13'b1110010001001,
13'b1110010010110,
13'b1110010010111,
13'b1110010011000,
13'b1110010011001,
13'b1110010011010,
13'b1110010100111,
13'b1110010101000,
13'b1110010101001,
13'b1110010101010,
13'b1110010111000,
13'b1110010111001,
13'b1111000100010,
13'b1111000100011,
13'b1111000100100,
13'b1111000100101,
13'b1111000110010,
13'b1111000110011,
13'b1111000110100,
13'b1111000110101,
13'b1111000110110,
13'b1111001000010,
13'b1111001000011,
13'b1111001000100,
13'b1111001000101,
13'b1111001000110,
13'b1111001000111,
13'b1111001010010,
13'b1111001010011,
13'b1111001010100,
13'b1111001010101,
13'b1111001010110,
13'b1111001010111,
13'b1111001100011,
13'b1111001100100,
13'b1111001100101,
13'b1111001100110,
13'b1111001100111,
13'b1111001101000,
13'b1111001110100,
13'b1111001110101,
13'b1111001110110,
13'b1111001110111,
13'b1111001111000,
13'b1111001111001,
13'b1111010000100,
13'b1111010000101,
13'b1111010000110,
13'b1111010000111,
13'b1111010001000,
13'b1111010001001,
13'b1111010010101,
13'b1111010010110,
13'b1111010010111,
13'b1111010011000,
13'b1111010011001,
13'b1111010100110,
13'b1111010100111,
13'b1111010101000,
13'b1111010101001,
13'b1111010111000,
13'b1111010111001: edge_mask_reg_512p3[269] <= 1'b1;
 		default: edge_mask_reg_512p3[269] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100111,
13'b11011101000,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100111,
13'b100011101000,
13'b101001000110,
13'b101001000111,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100111,
13'b101011101000,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110111,
13'b111010111000,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010001001,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010111000,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010001001,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110111,
13'b1001010111000,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010001001,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010110111,
13'b1010010111000,
13'b1011001110101,
13'b1011001110110,
13'b1011001110111,
13'b1011001111000,
13'b1011010000101,
13'b1011010000110,
13'b1011010000111,
13'b1011010001000,
13'b1011010001001,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010011001,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010110111,
13'b1011010111000,
13'b1011010111001,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100001110111,
13'b1100001111000,
13'b1100010000100,
13'b1100010000101,
13'b1100010000110,
13'b1100010000111,
13'b1100010001000,
13'b1100010001001,
13'b1100010010100,
13'b1100010010101,
13'b1100010010110,
13'b1100010010111,
13'b1100010011000,
13'b1100010011001,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010101001,
13'b1100010110111,
13'b1100010111000,
13'b1100010111001,
13'b1101001110100,
13'b1101001110101,
13'b1101001110110,
13'b1101001110111,
13'b1101001111000,
13'b1101010000100,
13'b1101010000101,
13'b1101010000110,
13'b1101010000111,
13'b1101010001000,
13'b1101010001001,
13'b1101010010100,
13'b1101010010101,
13'b1101010010110,
13'b1101010010111,
13'b1101010011000,
13'b1101010011001,
13'b1101010011010,
13'b1101010100100,
13'b1101010100101,
13'b1101010100110,
13'b1101010100111,
13'b1101010101000,
13'b1101010101001,
13'b1101010101010,
13'b1101010110111,
13'b1101010111000,
13'b1101010111001,
13'b1110001110100,
13'b1110001110101,
13'b1110001110110,
13'b1110001110111,
13'b1110001111000,
13'b1110010000011,
13'b1110010000100,
13'b1110010000101,
13'b1110010000110,
13'b1110010000111,
13'b1110010001000,
13'b1110010001001,
13'b1110010010011,
13'b1110010010100,
13'b1110010010101,
13'b1110010010110,
13'b1110010010111,
13'b1110010011000,
13'b1110010011001,
13'b1110010011010,
13'b1110010100100,
13'b1110010100101,
13'b1110010100110,
13'b1110010100111,
13'b1110010101000,
13'b1110010101001,
13'b1110010101010,
13'b1110010110111,
13'b1110010111000,
13'b1110010111001,
13'b1111001110100,
13'b1111001110101,
13'b1111001110110,
13'b1111001110111,
13'b1111001111000,
13'b1111010000011,
13'b1111010000100,
13'b1111010000101,
13'b1111010000110,
13'b1111010000111,
13'b1111010001000,
13'b1111010001001,
13'b1111010010011,
13'b1111010010100,
13'b1111010010101,
13'b1111010010110,
13'b1111010010111,
13'b1111010011000,
13'b1111010011001,
13'b1111010100011,
13'b1111010100100,
13'b1111010100101,
13'b1111010100110,
13'b1111010100111,
13'b1111010101000,
13'b1111010101001,
13'b1111010110111,
13'b1111010111000,
13'b1111010111001: edge_mask_reg_512p3[270] <= 1'b1;
 		default: edge_mask_reg_512p3[270] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b11001000000,
13'b11001000001,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010000,
13'b11001010001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100000,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b100000110000,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000000,
13'b100001000001,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010000,
13'b100001010001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100000,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010000,
13'b101001010001,
13'b101001010011,
13'b101001010100,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100000,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010111,
13'b111000011000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100111,
13'b111000101000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110111,
13'b111000111000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001010001,
13'b111001010010,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000001000001,
13'b1000001000010: edge_mask_reg_512p3[271] <= 1'b1;
 		default: edge_mask_reg_512p3[271] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[272] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000000,
13'b1010000001,
13'b1010000010,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010000,
13'b1010010001,
13'b1010010010,
13'b1010010011,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100000,
13'b1010100001,
13'b1010100010,
13'b1010100011,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110000,
13'b1010110001,
13'b1010110010,
13'b1010110011,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000000,
13'b1011000001,
13'b1011000010,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010000,
13'b1011010001,
13'b1011010010,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100000,
13'b1011100001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110000,
13'b10001110001,
13'b10001110010,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000000,
13'b10010000001,
13'b10010000010,
13'b10010000011,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010000,
13'b10010010001,
13'b10010010010,
13'b10010010011,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100000,
13'b10010100001,
13'b10010100010,
13'b10010100011,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110000,
13'b10010110001,
13'b10010110010,
13'b10010110011,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000000,
13'b10011000001,
13'b10011000010,
13'b10011000011,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010000,
13'b10011010001,
13'b10011010010,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100000,
13'b10011100001,
13'b10011100010,
13'b10011100011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110000,
13'b10011110001,
13'b10011110010,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100001,
13'b11001100010,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110000,
13'b11001110001,
13'b11001110010,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000000,
13'b11010000001,
13'b11010000010,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010000,
13'b11010010001,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100000,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110000,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000000,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010000,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100000,
13'b11011100001,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110000,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010001,
13'b100001010010,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100001,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110000,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000000,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010000,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100000,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110000,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000000,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110010,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000110,
13'b100100000111,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000000,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100001,
13'b101011100010,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000110,
13'b101100000111,
13'b110000110111,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110110,
13'b110011110111,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100111,
13'b111001101000,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110111,
13'b111001111000,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110001,
13'b111010110010,
13'b111010110110,
13'b111010110111,
13'b111011000110,
13'b111011000111,
13'b1000001010001,
13'b1000001010010,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010100001,
13'b1000010100010: edge_mask_reg_512p3[273] <= 1'b1;
 		default: edge_mask_reg_512p3[273] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10011101,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10101101,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b10111101,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100101000,
13'b100101001,
13'b100101010,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1001111101,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010001101,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010011101,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010101101,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1010111101,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b11001001010,
13'b11001001011,
13'b11001001100,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011010,
13'b100001011011,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001010,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011010,
13'b101010011011,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101010,
13'b101010101011,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111010,
13'b101010111011,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110101,
13'b101011111010,
13'b110001100101,
13'b110001100110,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110100,
13'b110011110101,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1001011000011,
13'b1001011010011: edge_mask_reg_512p3[274] <= 1'b1;
 		default: edge_mask_reg_512p3[274] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100000,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110000,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000000,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110110000101,
13'b110110000110,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111110010000,
13'b111110010001,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100101,
13'b111110100110,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1001110100000,
13'b1001110100001,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001111000000,
13'b1001111000001,
13'b1001111010000,
13'b1001111010001,
13'b1001111100000,
13'b1001111100001,
13'b1010110110000,
13'b1010110110001,
13'b1010111000000,
13'b1010111000001,
13'b1010111010000: edge_mask_reg_512p3[275] <= 1'b1;
 		default: edge_mask_reg_512p3[275] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10100000101,
13'b10100000110,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101100010101,
13'b101100010110,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111010101,
13'b110111010110,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000101,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010101,
13'b111101010110,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b1000100110000,
13'b1000100110001,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1001101000000,
13'b1001101000001,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001111000001,
13'b1010101010000,
13'b1010101010001,
13'b1010101100000,
13'b1010101100001,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1011101110000,
13'b1011101110001,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1100110000000,
13'b1100110010000,
13'b1100110010001,
13'b1100110100000,
13'b1100110100001,
13'b1100110100010,
13'b1100110110001,
13'b1101110010000,
13'b1101110100000: edge_mask_reg_512p3[276] <= 1'b1;
 		default: edge_mask_reg_512p3[276] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11010101,
13'b11010110,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010100,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011100101,
13'b1011100110,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100011110100,
13'b100011110101,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101011110101,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100000,
13'b110100100001,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111010101,
13'b110111010110,
13'b111100010001,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110101,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1001100100000,
13'b1001100100001,
13'b1001100110000,
13'b1001100110001,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001111000001,
13'b1010100110000,
13'b1010100110001,
13'b1010101000000,
13'b1010101000001,
13'b1010101010000,
13'b1010101010001,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1011101010000,
13'b1011101010001,
13'b1011101100000,
13'b1011101100001,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1100101110000,
13'b1100110000000,
13'b1100110000001,
13'b1100110010000,
13'b1100110010001,
13'b1100110100000,
13'b1100110100001,
13'b1100110100010,
13'b1100110110001,
13'b1101110000000,
13'b1101110010000,
13'b1101110100000: edge_mask_reg_512p3[277] <= 1'b1;
 		default: edge_mask_reg_512p3[277] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011001,
13'b10100011010,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010011,
13'b110011010100,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110101,
13'b1011010110110,
13'b1011011000101,
13'b1011011000110,
13'b1011011010101,
13'b1011011010110,
13'b1100001010101,
13'b1100001010110,
13'b1100001100101,
13'b1100001100110,
13'b1100001110101,
13'b1100001110110,
13'b1100010000101,
13'b1100010000110,
13'b1100010010101,
13'b1100010010110,
13'b1100010100101,
13'b1100010100110: edge_mask_reg_512p3[278] <= 1'b1;
 		default: edge_mask_reg_512p3[278] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100100,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110100,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000100,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100010101,
13'b1100010110,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100100100100,
13'b100100100101,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101100100101,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100101,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110101,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000101,
13'b111110000110,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010101,
13'b111110010110,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1001101010000,
13'b1001101010001,
13'b1001101100000,
13'b1001101100001,
13'b1001101110000,
13'b1001101110001,
13'b1001110000000,
13'b1001110000001,
13'b1001110010000,
13'b1001110010001,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001111000000,
13'b1001111000001,
13'b1001111010000,
13'b1001111010001,
13'b1001111100000,
13'b1001111100001,
13'b1010101100000,
13'b1010101110000,
13'b1010110000000,
13'b1010110010000,
13'b1010110100000,
13'b1010110100001,
13'b1010110110000,
13'b1010110110001,
13'b1010111000000,
13'b1010111000001,
13'b1010111010000: edge_mask_reg_512p3[279] <= 1'b1;
 		default: edge_mask_reg_512p3[279] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110001,
13'b11110010,
13'b11110011,
13'b11110100,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000001,
13'b100000010,
13'b100000011,
13'b100000100,
13'b100000111,
13'b100001000,
13'b100010001,
13'b100010010,
13'b100010011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100001,
13'b100100010,
13'b100100011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110001,
13'b100110010,
13'b100110011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010011,
13'b1011010100,
13'b1011010101,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100001,
13'b1011100010,
13'b1011100011,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110001,
13'b1011110010,
13'b1011110011,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000001,
13'b1100000010,
13'b1100000011,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010001,
13'b1100010010,
13'b1100010011,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100001,
13'b1100100010,
13'b1100100011,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110001,
13'b1100110010,
13'b1100110011,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000001,
13'b1101000010,
13'b1101000011,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000011,
13'b10011000100,
13'b10011000101,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100001,
13'b10011100010,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110001,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010001,
13'b10100010010,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100001,
13'b10100100010,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110001,
13'b10100110010,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010011,
13'b10101010100,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100001,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000001,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101001,
13'b11101101010,
13'b100010101000,
13'b100010101001,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000001,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101001,
13'b100101101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110011001000,
13'b110011001001,
13'b110011011001,
13'b110011100011,
13'b110011100100,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111001: edge_mask_reg_512p3[280] <= 1'b1;
 		default: edge_mask_reg_512p3[280] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110000,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000000,
13'b10011000001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010000,
13'b10011010001,
13'b10011010011,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100000,
13'b10011100001,
13'b10011100010,
13'b10011100011,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110000,
13'b10011110001,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000000,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110100,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000000,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010000,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100000,
13'b11011100001,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110000,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000000,
13'b11100000001,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010000,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110000,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000000,
13'b100100000001,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010000,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110000,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000000,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b111011010111,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100001000: edge_mask_reg_512p3[281] <= 1'b1;
 		default: edge_mask_reg_512p3[281] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[282] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[283] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001010,
13'b10110001011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001010,
13'b11110001011,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b101011001001,
13'b101011001010,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001000,
13'b110101001001,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100011001,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1010100011001,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1011011110011,
13'b1011011110100,
13'b1011011110101,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100001000,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1100011110011,
13'b1100011110100,
13'b1100100000011,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100010011,
13'b1100100010100,
13'b1100100010101,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1100100100011,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1101100000100,
13'b1101100000101,
13'b1101100000110,
13'b1101100010100,
13'b1101100010101,
13'b1101100010110,
13'b1101100010111,
13'b1101100100100,
13'b1101100100101,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100110110,
13'b1101100110111,
13'b1110100010101,
13'b1110100010110,
13'b1110100010111,
13'b1110100100101,
13'b1110100100110,
13'b1110100100111,
13'b1110100101000,
13'b1110100110110,
13'b1110100110111,
13'b1111100100111: edge_mask_reg_512p3[284] <= 1'b1;
 		default: edge_mask_reg_512p3[284] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011010,
13'b10001011011,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001010,
13'b10110001011,
13'b11001101010,
13'b11001101011,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111010,
13'b11101111011,
13'b11110001010,
13'b11110001011,
13'b100010001010,
13'b100010001011,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011010,
13'b100101011011,
13'b100101101010,
13'b100101101011,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b110010101001,
13'b110010101010,
13'b110010111001,
13'b110010111010,
13'b110010111011,
13'b110011001001,
13'b110011001010,
13'b110011001011,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001000,
13'b110101001001,
13'b111010101001,
13'b111010101010,
13'b111010111001,
13'b111010111010,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b1000010101000,
13'b1000010101001,
13'b1000010101010,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011011000,
13'b1000011011001,
13'b1000011011010,
13'b1000011101000,
13'b1000011101001,
13'b1000011101010,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000011111010,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100001010,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1001010101000,
13'b1001010101001,
13'b1001010101010,
13'b1001010111000,
13'b1001010111001,
13'b1001010111010,
13'b1001011001000,
13'b1001011001001,
13'b1001011001010,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011011010,
13'b1001011100111,
13'b1001011101000,
13'b1001011101001,
13'b1001011101010,
13'b1001011110111,
13'b1001011111000,
13'b1001011111001,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100010111,
13'b1001100011000,
13'b1001100011001,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1010010101000,
13'b1010010101001,
13'b1010010101010,
13'b1010010111000,
13'b1010010111001,
13'b1010010111010,
13'b1010011001000,
13'b1010011001001,
13'b1010011001010,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1010011011010,
13'b1010011100111,
13'b1010011101000,
13'b1010011101001,
13'b1010011110111,
13'b1010011111000,
13'b1010011111001,
13'b1010100000111,
13'b1010100001000,
13'b1010100001001,
13'b1010100010111,
13'b1010100011000,
13'b1010100011001,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100101001,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1011010101000,
13'b1011010101001,
13'b1011010101010,
13'b1011010111000,
13'b1011010111001,
13'b1011010111010,
13'b1011011001000,
13'b1011011001001,
13'b1011011001010,
13'b1011011010111,
13'b1011011011000,
13'b1011011011001,
13'b1011011011010,
13'b1011011100111,
13'b1011011101000,
13'b1011011101001,
13'b1011011110111,
13'b1011011111000,
13'b1011011111001,
13'b1011100000111,
13'b1011100001000,
13'b1011100001001,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100011001,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100101001,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000111,
13'b1011101001000,
13'b1100010101000,
13'b1100010101001,
13'b1100010111000,
13'b1100010111001,
13'b1100011000111,
13'b1100011001000,
13'b1100011001001,
13'b1100011010111,
13'b1100011011000,
13'b1100011011001,
13'b1100011100111,
13'b1100011101000,
13'b1100011101001,
13'b1100011110111,
13'b1100011111000,
13'b1100011111001,
13'b1100100000111,
13'b1100100001000,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1101010111000,
13'b1101010111001,
13'b1101011000111,
13'b1101011001000,
13'b1101011001001,
13'b1101011010111,
13'b1101011011000,
13'b1101011011001,
13'b1101011100111,
13'b1101011101000,
13'b1101011101001,
13'b1101011110111,
13'b1101011111000,
13'b1101011111001,
13'b1101100000110,
13'b1101100000111,
13'b1101100001000,
13'b1101100010110,
13'b1101100010111,
13'b1101100011000,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100110110,
13'b1101100110111,
13'b1110010110111,
13'b1110010111000,
13'b1110010111001,
13'b1110011000111,
13'b1110011001000,
13'b1110011001001,
13'b1110011010111,
13'b1110011011000,
13'b1110011011001,
13'b1110011100111,
13'b1110011101000,
13'b1110011110111,
13'b1110011111000,
13'b1110100000110,
13'b1110100000111,
13'b1110100001000,
13'b1110100010110,
13'b1110100010111,
13'b1110100011000,
13'b1110100100110,
13'b1110100100111,
13'b1110100101000,
13'b1110100110110,
13'b1110100110111,
13'b1111010111000,
13'b1111010111001,
13'b1111011000111,
13'b1111011001000,
13'b1111011001001,
13'b1111011010111,
13'b1111011011000,
13'b1111011011001,
13'b1111011100111,
13'b1111011101000,
13'b1111011110111,
13'b1111011111000,
13'b1111100000111,
13'b1111100001000,
13'b1111100010111,
13'b1111100011000,
13'b1111100100111,
13'b1111100101000: edge_mask_reg_512p3[285] <= 1'b1;
 		default: edge_mask_reg_512p3[285] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b110000100110: edge_mask_reg_512p3[286] <= 1'b1;
 		default: edge_mask_reg_512p3[286] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101101001,
13'b101101010,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11110001010,
13'b11110001011,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111011001,
13'b101111011010,
13'b101111011011,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b110111011011,
13'b111111001001,
13'b111111001010,
13'b111111001011,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111011011,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b111111101010,
13'b111111101011,
13'b1000111001001,
13'b1000111001010,
13'b1000111001011,
13'b1000111011000,
13'b1000111011001,
13'b1000111011010,
13'b1000111011011,
13'b1000111100111,
13'b1000111101000,
13'b1000111101001,
13'b1000111101010,
13'b1000111101011,
13'b1001111001001,
13'b1001111001010,
13'b1001111001011,
13'b1001111011000,
13'b1001111011001,
13'b1001111011010,
13'b1001111011011,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1001111101001,
13'b1001111101010,
13'b1001111101011,
13'b1010111001000,
13'b1010111001001,
13'b1010111001010,
13'b1010111001011,
13'b1010111010111,
13'b1010111011000,
13'b1010111011001,
13'b1010111011010,
13'b1010111011011,
13'b1010111100110,
13'b1010111100111,
13'b1010111101000,
13'b1010111101001,
13'b1010111101010,
13'b1010111101011,
13'b1010111110110,
13'b1010111110111,
13'b1010111111000,
13'b1010111111001,
13'b1010111111010,
13'b1010111111011,
13'b1011111001000,
13'b1011111001001,
13'b1011111001010,
13'b1011111001011,
13'b1011111010111,
13'b1011111011000,
13'b1011111011001,
13'b1011111011010,
13'b1011111011011,
13'b1011111100110,
13'b1011111100111,
13'b1011111101000,
13'b1011111101001,
13'b1011111101010,
13'b1011111101011,
13'b1011111110101,
13'b1011111110110,
13'b1011111110111,
13'b1011111111000,
13'b1011111111001,
13'b1011111111010,
13'b1011111111011,
13'b1100111001000,
13'b1100111001001,
13'b1100111001010,
13'b1100111001011,
13'b1100111010111,
13'b1100111011000,
13'b1100111011001,
13'b1100111011010,
13'b1100111011011,
13'b1100111100110,
13'b1100111100111,
13'b1100111101000,
13'b1100111101001,
13'b1100111101010,
13'b1100111101011,
13'b1100111110101,
13'b1100111110110,
13'b1100111110111,
13'b1100111111000,
13'b1100111111001,
13'b1100111111010,
13'b1100111111011,
13'b1101111001001,
13'b1101111001010,
13'b1101111011000,
13'b1101111011001,
13'b1101111011010,
13'b1101111011011,
13'b1101111100110,
13'b1101111100111,
13'b1101111101000,
13'b1101111101001,
13'b1101111101010,
13'b1101111101011,
13'b1101111110101,
13'b1101111110110,
13'b1101111110111,
13'b1101111111000,
13'b1101111111001,
13'b1101111111010,
13'b1101111111011,
13'b1110111011000,
13'b1110111011001,
13'b1110111011010,
13'b1110111100110,
13'b1110111100111,
13'b1110111101000,
13'b1110111101001,
13'b1110111101010,
13'b1110111110101,
13'b1110111110110,
13'b1110111110111,
13'b1110111111000,
13'b1110111111001,
13'b1111111011000,
13'b1111111011001,
13'b1111111100110,
13'b1111111100111,
13'b1111111101000,
13'b1111111101001,
13'b1111111101010,
13'b1111111110101,
13'b1111111110110,
13'b1111111110111,
13'b1111111111000,
13'b1111111111001: edge_mask_reg_512p3[287] <= 1'b1;
 		default: edge_mask_reg_512p3[287] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100110111100,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b100111001100,
13'b101101011001,
13'b101101011010,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111011001,
13'b101111011010,
13'b101111011011,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111001011,
13'b110111011001,
13'b110111011010,
13'b110111011011,
13'b111101110111,
13'b111101111000,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110111000,
13'b111110111001,
13'b111110111010,
13'b111111001000,
13'b111111001001,
13'b111111001010,
13'b111111001011,
13'b111111011000,
13'b111111011001,
13'b111111011010,
13'b111111011011,
13'b111111101001,
13'b111111101010,
13'b111111101011,
13'b1000101110111,
13'b1000101111000,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110011001,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110101010,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000110111010,
13'b1000111001000,
13'b1000111001001,
13'b1000111001010,
13'b1000111001011,
13'b1000111011000,
13'b1000111011001,
13'b1000111011010,
13'b1000111011011,
13'b1000111101001,
13'b1000111101010,
13'b1000111101011,
13'b1001101110111,
13'b1001101111000,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110001001,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110011001,
13'b1001110100111,
13'b1001110101000,
13'b1001110101001,
13'b1001110101010,
13'b1001110110111,
13'b1001110111000,
13'b1001110111001,
13'b1001110111010,
13'b1001111001000,
13'b1001111001001,
13'b1001111001010,
13'b1001111001011,
13'b1001111011000,
13'b1001111011001,
13'b1001111011010,
13'b1001111011011,
13'b1001111101001,
13'b1001111101010,
13'b1001111101011,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1010110011001,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110101001,
13'b1010110101010,
13'b1010110110111,
13'b1010110111000,
13'b1010110111001,
13'b1010110111010,
13'b1010111000111,
13'b1010111001000,
13'b1010111001001,
13'b1010111001010,
13'b1010111001011,
13'b1010111011000,
13'b1010111011001,
13'b1010111011010,
13'b1010111011011,
13'b1010111101001,
13'b1010111101010,
13'b1010111101011,
13'b1010111111001,
13'b1010111111010,
13'b1010111111011,
13'b1011101110110,
13'b1011101110111,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1011110011001,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110101001,
13'b1011110110110,
13'b1011110110111,
13'b1011110111000,
13'b1011110111001,
13'b1011110111010,
13'b1011111000111,
13'b1011111001000,
13'b1011111001001,
13'b1011111001010,
13'b1011111001011,
13'b1011111011000,
13'b1011111011001,
13'b1011111011010,
13'b1011111011011,
13'b1011111101000,
13'b1011111101001,
13'b1011111101010,
13'b1011111101011,
13'b1011111111001,
13'b1011111111010,
13'b1011111111011,
13'b1100101110110,
13'b1100101110111,
13'b1100110000101,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1100110100101,
13'b1100110100110,
13'b1100110100111,
13'b1100110101000,
13'b1100110101001,
13'b1100110110110,
13'b1100110110111,
13'b1100110111000,
13'b1100110111001,
13'b1100110111010,
13'b1100111000111,
13'b1100111001000,
13'b1100111001001,
13'b1100111001010,
13'b1100111001011,
13'b1100111011000,
13'b1100111011001,
13'b1100111011010,
13'b1100111011011,
13'b1100111101000,
13'b1100111101001,
13'b1100111101010,
13'b1100111101011,
13'b1100111111001,
13'b1100111111010,
13'b1100111111011,
13'b1101110000101,
13'b1101110000110,
13'b1101110000111,
13'b1101110010100,
13'b1101110010101,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1101110100111,
13'b1101110101000,
13'b1101110101001,
13'b1101110110101,
13'b1101110110110,
13'b1101110110111,
13'b1101110111000,
13'b1101110111001,
13'b1101110111010,
13'b1101111000110,
13'b1101111000111,
13'b1101111001000,
13'b1101111001001,
13'b1101111001010,
13'b1101111010111,
13'b1101111011000,
13'b1101111011001,
13'b1101111011010,
13'b1101111011011,
13'b1101111101000,
13'b1101111101001,
13'b1101111101010,
13'b1101111101011,
13'b1101111111001,
13'b1101111111010,
13'b1101111111011,
13'b1110110000101,
13'b1110110000110,
13'b1110110010100,
13'b1110110010101,
13'b1110110010110,
13'b1110110010111,
13'b1110110100100,
13'b1110110100101,
13'b1110110100110,
13'b1110110100111,
13'b1110110101000,
13'b1110110110101,
13'b1110110110110,
13'b1110110110111,
13'b1110110111000,
13'b1110110111001,
13'b1110111000110,
13'b1110111000111,
13'b1110111001000,
13'b1110111001001,
13'b1110111010111,
13'b1110111011000,
13'b1110111011001,
13'b1110111011010,
13'b1110111101000,
13'b1110111101001,
13'b1110111101010,
13'b1110111111000,
13'b1110111111001,
13'b1111110000101,
13'b1111110010101,
13'b1111110010110,
13'b1111110010111,
13'b1111110100101,
13'b1111110100110,
13'b1111110100111,
13'b1111110110101,
13'b1111110110110,
13'b1111110110111,
13'b1111110111000,
13'b1111111000110,
13'b1111111000111,
13'b1111111001000,
13'b1111111001001,
13'b1111111010111,
13'b1111111011000,
13'b1111111011001,
13'b1111111100111,
13'b1111111101000,
13'b1111111101001,
13'b1111111101010,
13'b1111111111000,
13'b1111111111001: edge_mask_reg_512p3[288] <= 1'b1;
 		default: edge_mask_reg_512p3[288] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[289] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110101000,
13'b11110101001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110101000,
13'b100110101001,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110011000,
13'b101110011001,
13'b110011010111,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110001000,
13'b110110001001,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b1000100000110,
13'b1000100000111,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110111,
13'b1010101111000,
13'b1011011110110,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101011001,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010100,
13'b1100100010101,
13'b1100100010110,
13'b1100100010111,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101011001,
13'b1100101100111,
13'b1100101101000,
13'b1100101101001,
13'b1100101110111,
13'b1100101111000,
13'b1101100000100,
13'b1101100000101,
13'b1101100000110,
13'b1101100010100,
13'b1101100010101,
13'b1101100010110,
13'b1101100010111,
13'b1101100100100,
13'b1101100100101,
13'b1101100100110,
13'b1101100100111,
13'b1101100110100,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101011001,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101101001,
13'b1101101110111,
13'b1101101111000,
13'b1110100000100,
13'b1110100000101,
13'b1110100000110,
13'b1110100010100,
13'b1110100010101,
13'b1110100010110,
13'b1110100010111,
13'b1110100100100,
13'b1110100100101,
13'b1110100100110,
13'b1110100100111,
13'b1110100110100,
13'b1110100110101,
13'b1110100110110,
13'b1110100110111,
13'b1110100111000,
13'b1110101000101,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101011001,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110111,
13'b1111100000100,
13'b1111100000101,
13'b1111100010011,
13'b1111100010100,
13'b1111100010101,
13'b1111100010110,
13'b1111100100011,
13'b1111100100100,
13'b1111100100101,
13'b1111100100110,
13'b1111100100111,
13'b1111100110100,
13'b1111100110101,
13'b1111100110110,
13'b1111100110111,
13'b1111100111000,
13'b1111101000101,
13'b1111101000110,
13'b1111101000111,
13'b1111101001000,
13'b1111101010110,
13'b1111101010111,
13'b1111101011000,
13'b1111101100111,
13'b1111101101000: edge_mask_reg_512p3[290] <= 1'b1;
 		default: edge_mask_reg_512p3[290] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[291] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101101000,
13'b101101001,
13'b1101111000,
13'b1101111001,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b101111011011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110110100,
13'b1001110110101,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1011111110111,
13'b1100111010011,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110,
13'b1101111100011,
13'b1101111100100,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1101111110110,
13'b1110111110100,
13'b1110111110101: edge_mask_reg_512p3[292] <= 1'b1;
 		default: edge_mask_reg_512p3[292] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100000,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110000,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110110,
13'b100011110111,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100110,
13'b110011100111,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010000,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100000,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010110000,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000011000001,
13'b1000011000010,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001010000000,
13'b1001010000001,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010010001,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010110001,
13'b1001010110010,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001110000,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010010010,
13'b1010010010011,
13'b1011000110011,
13'b1011001000010,
13'b1011001000011,
13'b1011001010000,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001100000,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001110010,
13'b1011001110011: edge_mask_reg_512p3[293] <= 1'b1;
 		default: edge_mask_reg_512p3[293] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110000,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000000,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010000,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100000,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110000,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110110,
13'b100011110111,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b110000110111,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100110,
13'b110011100111,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100111,
13'b111001101000,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110111,
13'b111001111000,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000111,
13'b111010001000,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b1000001010001,
13'b1000001010010,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010010000,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010100000,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010110000,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000011000001,
13'b1000011000010: edge_mask_reg_512p3[294] <= 1'b1;
 		default: edge_mask_reg_512p3[294] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[295] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011010,
13'b10101011011,
13'b10101101010,
13'b10101101011,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100111,
13'b101100101000,
13'b110010100110,
13'b110010100111,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100100,
13'b110100100101,
13'b110100100111,
13'b110100101000,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1001010100100,
13'b1001010100101,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100110,
13'b1010010110100,
13'b1010010110101,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110101,
13'b1010011110110,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1011011000101,
13'b1011011010101,
13'b1011011100101: edge_mask_reg_512p3[296] <= 1'b1;
 		default: edge_mask_reg_512p3[296] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101010,
13'b1101101011,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011010,
13'b10101011011,
13'b10101101010,
13'b10101101011,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011010,
13'b11101011011,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001010,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100100,
13'b101100100111,
13'b101100101000,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110011,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000011,
13'b110011000100,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010011,
13'b110011010100,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100100,
13'b110100100101,
13'b110100100111,
13'b110100101000,
13'b111010010110,
13'b111010010111,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b1000010010110,
13'b1000010010111,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100110,
13'b1000100100111,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100110,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010110,
13'b1010100010111,
13'b1011010100101,
13'b1011010100110,
13'b1011010110101,
13'b1011010110110,
13'b1011011000101,
13'b1011011000110,
13'b1011011010101,
13'b1011011010110,
13'b1011011100101,
13'b1011011100110,
13'b1011011110101,
13'b1011011110110: edge_mask_reg_512p3[297] <= 1'b1;
 		default: edge_mask_reg_512p3[297] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11010101,
13'b11010110,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010100,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100100,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110100,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000100,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011100101,
13'b1011100110,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000011,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110010011,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110100011,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b100011110100,
13'b100011110101,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b101011110101,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101111000100,
13'b101111000101,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100100000,
13'b110100100001,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110100001,
13'b110110100010,
13'b110110100100,
13'b110110100101,
13'b110110110100,
13'b110110110101,
13'b111100010001,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110101,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000101,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010101,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110100000,
13'b1000110100001,
13'b1001100100000,
13'b1001100100001,
13'b1001100110000,
13'b1001100110001,
13'b1001101000000,
13'b1001101000001,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110100000,
13'b1010100110000,
13'b1010101000000,
13'b1010101000001,
13'b1010101010000,
13'b1010101010001,
13'b1010101100000,
13'b1010101100001,
13'b1010101110000,
13'b1010101110001,
13'b1010110000000,
13'b1010110000001,
13'b1010110010000,
13'b1010110010001: edge_mask_reg_512p3[298] <= 1'b1;
 		default: edge_mask_reg_512p3[298] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110111000,
13'b100011101000,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b101011101000,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110101000,
13'b101110101001,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110011000,
13'b110110011001,
13'b111100011000,
13'b111100011001,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b1000100101000,
13'b1000100101001,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101001011,
13'b1000101011000,
13'b1000101011001,
13'b1000101011010,
13'b1000101011011,
13'b1000101101000,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1001100011001,
13'b1001100101000,
13'b1001100101001,
13'b1001100101010,
13'b1001100111000,
13'b1001100111001,
13'b1001100111010,
13'b1001101001000,
13'b1001101001001,
13'b1001101001010,
13'b1001101001011,
13'b1001101011000,
13'b1001101011001,
13'b1001101011010,
13'b1001101011011,
13'b1001101101001,
13'b1001101101010,
13'b1001101101011,
13'b1001101111001,
13'b1001101111010,
13'b1001101111011,
13'b1010100011001,
13'b1010100101000,
13'b1010100101001,
13'b1010100101010,
13'b1010100111000,
13'b1010100111001,
13'b1010100111010,
13'b1010100111011,
13'b1010101001000,
13'b1010101001001,
13'b1010101001010,
13'b1010101001011,
13'b1010101011000,
13'b1010101011001,
13'b1010101011010,
13'b1010101011011,
13'b1010101101001,
13'b1010101101010,
13'b1010101101011,
13'b1010101101100,
13'b1010101111001,
13'b1010101111010,
13'b1010101111011,
13'b1010101111100,
13'b1011100011000,
13'b1011100011001,
13'b1011100101000,
13'b1011100101001,
13'b1011100101010,
13'b1011100111000,
13'b1011100111001,
13'b1011100111010,
13'b1011100111011,
13'b1011101001000,
13'b1011101001001,
13'b1011101001010,
13'b1011101001011,
13'b1011101001100,
13'b1011101011000,
13'b1011101011001,
13'b1011101011010,
13'b1011101011011,
13'b1011101011100,
13'b1011101101001,
13'b1011101101010,
13'b1011101101011,
13'b1011101101100,
13'b1011101111010,
13'b1011101111011,
13'b1011101111100,
13'b1100100011000,
13'b1100100011001,
13'b1100100101000,
13'b1100100101001,
13'b1100100101010,
13'b1100100111000,
13'b1100100111001,
13'b1100100111010,
13'b1100100111011,
13'b1100101001000,
13'b1100101001001,
13'b1100101001010,
13'b1100101001011,
13'b1100101001100,
13'b1100101011000,
13'b1100101011001,
13'b1100101011010,
13'b1100101011011,
13'b1100101011100,
13'b1100101101001,
13'b1100101101010,
13'b1100101101011,
13'b1100101101100,
13'b1100101111010,
13'b1100101111011,
13'b1100101111100,
13'b1101100011001,
13'b1101100101000,
13'b1101100101001,
13'b1101100101010,
13'b1101100111000,
13'b1101100111001,
13'b1101100111010,
13'b1101100111011,
13'b1101101001000,
13'b1101101001001,
13'b1101101001010,
13'b1101101001011,
13'b1101101001100,
13'b1101101011001,
13'b1101101011010,
13'b1101101011011,
13'b1101101011100,
13'b1101101101001,
13'b1101101101010,
13'b1101101101011,
13'b1101101101100,
13'b1101101111010,
13'b1101101111011,
13'b1101101111100,
13'b1110100011001,
13'b1110100101000,
13'b1110100101001,
13'b1110100101010,
13'b1110100110111,
13'b1110100111000,
13'b1110100111001,
13'b1110100111010,
13'b1110100111011,
13'b1110101000111,
13'b1110101001000,
13'b1110101001001,
13'b1110101001010,
13'b1110101001011,
13'b1110101011000,
13'b1110101011001,
13'b1110101011010,
13'b1110101011011,
13'b1110101011100,
13'b1110101101001,
13'b1110101101010,
13'b1110101101011,
13'b1110101101100,
13'b1110101111010,
13'b1110101111011,
13'b1111100101000,
13'b1111100101001,
13'b1111100101010,
13'b1111100110111,
13'b1111100111000,
13'b1111100111001,
13'b1111100111010,
13'b1111101000111,
13'b1111101001000,
13'b1111101001001,
13'b1111101001010,
13'b1111101001011,
13'b1111101011000,
13'b1111101011001,
13'b1111101011010,
13'b1111101011011,
13'b1111101101001,
13'b1111101101010,
13'b1111101101011,
13'b1111101111010,
13'b1111101111011: edge_mask_reg_512p3[299] <= 1'b1;
 		default: edge_mask_reg_512p3[299] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010100111,
13'b1010101000,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110111000,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b101010111000,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110101000,
13'b101110101001,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110011000,
13'b110110011001,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b1000011101001,
13'b1000011101010,
13'b1000011111000,
13'b1000011111001,
13'b1000011111010,
13'b1000100001000,
13'b1000100001001,
13'b1000100001010,
13'b1000100011000,
13'b1000100011001,
13'b1000100011010,
13'b1000100101000,
13'b1000100101001,
13'b1000100101010,
13'b1000100101011,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000100111011,
13'b1000101001001,
13'b1000101001010,
13'b1000101001011,
13'b1000101011001,
13'b1000101011010,
13'b1000101011011,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1001011101001,
13'b1001011101010,
13'b1001011111000,
13'b1001011111001,
13'b1001011111010,
13'b1001100001000,
13'b1001100001001,
13'b1001100001010,
13'b1001100001011,
13'b1001100011001,
13'b1001100011010,
13'b1001100011011,
13'b1001100101001,
13'b1001100101010,
13'b1001100101011,
13'b1001100111001,
13'b1001100111010,
13'b1001100111011,
13'b1001101001001,
13'b1001101001010,
13'b1001101001011,
13'b1001101011001,
13'b1001101011010,
13'b1001101011011,
13'b1001101101001,
13'b1001101101010,
13'b1001101101011,
13'b1001101111001,
13'b1001101111010,
13'b1001101111011,
13'b1010011101001,
13'b1010011101010,
13'b1010011101011,
13'b1010011111001,
13'b1010011111010,
13'b1010011111011,
13'b1010100001001,
13'b1010100001010,
13'b1010100001011,
13'b1010100011001,
13'b1010100011010,
13'b1010100011011,
13'b1010100101001,
13'b1010100101010,
13'b1010100101011,
13'b1010100111001,
13'b1010100111010,
13'b1010100111011,
13'b1010101001001,
13'b1010101001010,
13'b1010101001011,
13'b1010101011001,
13'b1010101011010,
13'b1010101011011,
13'b1010101101001,
13'b1010101101010,
13'b1010101101011,
13'b1010101101100,
13'b1010101111010,
13'b1010101111011,
13'b1010101111100,
13'b1011011101001,
13'b1011011101010,
13'b1011011101011,
13'b1011011111001,
13'b1011011111010,
13'b1011011111011,
13'b1011100001001,
13'b1011100001010,
13'b1011100001011,
13'b1011100011001,
13'b1011100011010,
13'b1011100011011,
13'b1011100101001,
13'b1011100101010,
13'b1011100101011,
13'b1011100101100,
13'b1011100111001,
13'b1011100111010,
13'b1011100111011,
13'b1011100111100,
13'b1011101001001,
13'b1011101001010,
13'b1011101001011,
13'b1011101001100,
13'b1011101011001,
13'b1011101011010,
13'b1011101011011,
13'b1011101011100,
13'b1011101101010,
13'b1011101101011,
13'b1011101101100,
13'b1011101111010,
13'b1011101111011,
13'b1011101111100,
13'b1100011101001,
13'b1100011101010,
13'b1100011101011,
13'b1100011111001,
13'b1100011111010,
13'b1100011111011,
13'b1100100001001,
13'b1100100001010,
13'b1100100001011,
13'b1100100001100,
13'b1100100011001,
13'b1100100011010,
13'b1100100011011,
13'b1100100011100,
13'b1100100101001,
13'b1100100101010,
13'b1100100101011,
13'b1100100101100,
13'b1100100111010,
13'b1100100111011,
13'b1100100111100,
13'b1100101001010,
13'b1100101001011,
13'b1100101001100,
13'b1100101011010,
13'b1100101011011,
13'b1100101011100,
13'b1100101101010,
13'b1100101101011,
13'b1100101101100,
13'b1100101111010,
13'b1100101111011,
13'b1100101111100,
13'b1101011101001,
13'b1101011101010,
13'b1101011101011,
13'b1101011111001,
13'b1101011111010,
13'b1101011111011,
13'b1101100001001,
13'b1101100001010,
13'b1101100001011,
13'b1101100001100,
13'b1101100011001,
13'b1101100011010,
13'b1101100011011,
13'b1101100011100,
13'b1101100101001,
13'b1101100101010,
13'b1101100101011,
13'b1101100101100,
13'b1101100111010,
13'b1101100111011,
13'b1101100111100,
13'b1101101001010,
13'b1101101001011,
13'b1101101001100,
13'b1101101011010,
13'b1101101011011,
13'b1101101011100,
13'b1101101101010,
13'b1101101101011,
13'b1101101101100,
13'b1101101111010,
13'b1101101111011,
13'b1101101111100,
13'b1110011101010,
13'b1110011101011,
13'b1110011111001,
13'b1110011111010,
13'b1110011111011,
13'b1110100001001,
13'b1110100001010,
13'b1110100001011,
13'b1110100011001,
13'b1110100011010,
13'b1110100011011,
13'b1110100101001,
13'b1110100101010,
13'b1110100101011,
13'b1110100101100,
13'b1110100111001,
13'b1110100111010,
13'b1110100111011,
13'b1110100111100,
13'b1110101001001,
13'b1110101001010,
13'b1110101001011,
13'b1110101001100,
13'b1110101011001,
13'b1110101011010,
13'b1110101011011,
13'b1110101011100,
13'b1110101101010,
13'b1110101101011,
13'b1110101101100,
13'b1110101111010,
13'b1110101111011,
13'b1111011111001,
13'b1111011111010,
13'b1111100001000,
13'b1111100001001,
13'b1111100001010,
13'b1111100001011,
13'b1111100011000,
13'b1111100011001,
13'b1111100011010,
13'b1111100011011,
13'b1111100101000,
13'b1111100101001,
13'b1111100101010,
13'b1111100101011,
13'b1111100111001,
13'b1111100111010,
13'b1111100111011,
13'b1111101001001,
13'b1111101001010,
13'b1111101001011,
13'b1111101011001,
13'b1111101011010,
13'b1111101011011,
13'b1111101101001,
13'b1111101101010,
13'b1111101101011,
13'b1111101111010,
13'b1111101111011: edge_mask_reg_512p3[300] <= 1'b1;
 		default: edge_mask_reg_512p3[300] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110011000,
13'b110110011001,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b1000100111010,
13'b1000100111011,
13'b1000101001001,
13'b1000101001010,
13'b1000101001011,
13'b1000101011001,
13'b1000101011010,
13'b1000101011011,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1001100111010,
13'b1001100111011,
13'b1001101001001,
13'b1001101001010,
13'b1001101001011,
13'b1001101001100,
13'b1001101011001,
13'b1001101011010,
13'b1001101011011,
13'b1001101011100,
13'b1001101101001,
13'b1001101101010,
13'b1001101101011,
13'b1001101101100,
13'b1001101111001,
13'b1001101111010,
13'b1001101111011,
13'b1010100111010,
13'b1010100111011,
13'b1010100111100,
13'b1010101001001,
13'b1010101001010,
13'b1010101001011,
13'b1010101001100,
13'b1010101011001,
13'b1010101011010,
13'b1010101011011,
13'b1010101011100,
13'b1010101101001,
13'b1010101101010,
13'b1010101101011,
13'b1010101101100,
13'b1010101111010,
13'b1010101111011,
13'b1010101111100,
13'b1011100111010,
13'b1011100111011,
13'b1011100111100,
13'b1011101001001,
13'b1011101001010,
13'b1011101001011,
13'b1011101001100,
13'b1011101011001,
13'b1011101011010,
13'b1011101011011,
13'b1011101011100,
13'b1011101011101,
13'b1011101101010,
13'b1011101101011,
13'b1011101101100,
13'b1011101101101,
13'b1011101111010,
13'b1011101111011,
13'b1011101111100,
13'b1100100111011,
13'b1100100111100,
13'b1100101001010,
13'b1100101001011,
13'b1100101001100,
13'b1100101011010,
13'b1100101011011,
13'b1100101011100,
13'b1100101011101,
13'b1100101101010,
13'b1100101101011,
13'b1100101101100,
13'b1100101101101,
13'b1100101111010,
13'b1100101111011,
13'b1100101111100,
13'b1101100111011,
13'b1101100111100,
13'b1101101001010,
13'b1101101001011,
13'b1101101001100,
13'b1101101011010,
13'b1101101011011,
13'b1101101011100,
13'b1101101101010,
13'b1101101101011,
13'b1101101101100,
13'b1101101111010,
13'b1101101111011,
13'b1101101111100,
13'b1110101001010,
13'b1110101001011,
13'b1110101001100,
13'b1110101011010,
13'b1110101011011,
13'b1110101011100,
13'b1110101101010,
13'b1110101101011,
13'b1110101101100,
13'b1110101111010,
13'b1110101111011,
13'b1111101001010,
13'b1111101001011,
13'b1111101011010,
13'b1111101011011,
13'b1111101011100,
13'b1111101101001,
13'b1111101101010,
13'b1111101101011,
13'b1111101101100,
13'b1111101111010,
13'b1111101111011: edge_mask_reg_512p3[301] <= 1'b1;
 		default: edge_mask_reg_512p3[301] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000110,
13'b1101000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b100001010110,
13'b100001010111,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b101001010110,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110110,
13'b110100110111,
13'b111001110010,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b1000001110010,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010010000,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010100000,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110000,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1001010000000,
13'b1001010000001,
13'b1001010000010,
13'b1001010000011,
13'b1001010010000,
13'b1001010010001,
13'b1001010010010,
13'b1001010010011,
13'b1001010100000,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010110000,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1010010000001,
13'b1010010000010,
13'b1010010010000,
13'b1010010010001,
13'b1010010010010,
13'b1010010100000,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010110000,
13'b1010010110001,
13'b1010010110010,
13'b1010010110011,
13'b1010011000000,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1011010010000,
13'b1011010010001,
13'b1011010010010,
13'b1011010100000,
13'b1011010100001,
13'b1011010100010,
13'b1011010110000,
13'b1011010110001,
13'b1011010110010,
13'b1011010110011,
13'b1011011000000,
13'b1011011000001,
13'b1011011000010,
13'b1011011000011,
13'b1011011010000,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1100010100000,
13'b1100010100001,
13'b1100010110000,
13'b1100010110001,
13'b1100010110010,
13'b1100011000000,
13'b1100011000001,
13'b1100011000010,
13'b1100011000011,
13'b1100011010000,
13'b1100011010001,
13'b1100011010010,
13'b1100011010011,
13'b1100011100000,
13'b1100011100001,
13'b1100011100010,
13'b1100011100011,
13'b1100011110000,
13'b1100011110001,
13'b1100011110010,
13'b1100011110011,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1101010100000,
13'b1101010110000,
13'b1101010110001,
13'b1101011000000,
13'b1101011000001,
13'b1101011010000,
13'b1101011010001,
13'b1101011010010,
13'b1101011100000,
13'b1101011100001,
13'b1101011100010,
13'b1101011100011,
13'b1101011110000,
13'b1101011110001,
13'b1101011110010,
13'b1101011110011,
13'b1101100000010,
13'b1101100000011,
13'b1110011000000,
13'b1110011000001,
13'b1110011010000,
13'b1110011010001,
13'b1110011010010,
13'b1110011100000,
13'b1110011100001,
13'b1110011100010,
13'b1110011110000,
13'b1110011110001,
13'b1110011110010,
13'b1111011010000,
13'b1111011010001,
13'b1111011100000,
13'b1111011100001,
13'b1111011110000,
13'b1111011110001: edge_mask_reg_512p3[302] <= 1'b1;
 		default: edge_mask_reg_512p3[302] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b100001010110,
13'b100001010111,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b101001010110,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010110,
13'b101100010111,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110011,
13'b110011110100,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010110,
13'b110100010111,
13'b111001110010,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b1000001110010,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010010000,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010100000,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010110000,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000000,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010000,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1001010000000,
13'b1001010000001,
13'b1001010000010,
13'b1001010000011,
13'b1001010010000,
13'b1001010010001,
13'b1001010010010,
13'b1001010010011,
13'b1001010100000,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010110000,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011110001,
13'b1001011110010,
13'b1010010000001,
13'b1010010000010,
13'b1010010010000,
13'b1010010010001,
13'b1010010010010,
13'b1010010100000,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010110000,
13'b1010010110001,
13'b1010010110010,
13'b1010010110011,
13'b1010011000000,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011110001,
13'b1011010010000,
13'b1011010010001,
13'b1011010100000,
13'b1011010100001,
13'b1011010100010,
13'b1011010110000,
13'b1011010110001,
13'b1011010110010,
13'b1011011000000,
13'b1011011000001,
13'b1011011000010,
13'b1011011010000,
13'b1011011010001,
13'b1100010100000: edge_mask_reg_512p3[303] <= 1'b1;
 		default: edge_mask_reg_512p3[303] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000110,
13'b1010000111,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110110,
13'b1011110111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b110001010110,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011100110,
13'b110011100111,
13'b111001110010,
13'b111001110011,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000010,
13'b111011000011,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010010000,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010100000,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010110000,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001010000000,
13'b1001010000001,
13'b1001010000010,
13'b1001010000011,
13'b1001010010000,
13'b1001010010001,
13'b1001010010010,
13'b1001010010011,
13'b1001010100000,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010110000,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001011000001,
13'b1001011000010,
13'b1010001110001,
13'b1010001110010,
13'b1010010000000,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010010000,
13'b1010010010001,
13'b1010010010010,
13'b1010010100000,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010110000,
13'b1010010110001,
13'b1010010110010,
13'b1010010110011,
13'b1010011000001,
13'b1011001110001,
13'b1011001110010,
13'b1011010000000,
13'b1011010000001,
13'b1011010000010,
13'b1011010010000,
13'b1011010010001,
13'b1011010010010,
13'b1011010100000,
13'b1011010100001,
13'b1011010100010,
13'b1011010110000,
13'b1011010110001,
13'b1011010110010,
13'b1100010000000,
13'b1100010000001,
13'b1100010010000,
13'b1100010010001,
13'b1100010100000,
13'b1100010100001,
13'b1101010000000,
13'b1101010010000,
13'b1101010100000: edge_mask_reg_512p3[304] <= 1'b1;
 		default: edge_mask_reg_512p3[304] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[305] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111000,
13'b100110111001,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b110011010111,
13'b110011011000,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110011000,
13'b110110011001,
13'b111011010111,
13'b111011011000,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000101,
13'b111110000110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1001011010110,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000100,
13'b1001110000101,
13'b1010011010110,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000010,
13'b1010110000100,
13'b1010110000101,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000011,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010011,
13'b1100100010100,
13'b1100100010101,
13'b1100100010110,
13'b1100100010111,
13'b1100100100011,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100110011,
13'b1100100110100,
13'b1100100110101,
13'b1100100110110,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110010,
13'b1100101110100,
13'b1100101110101,
13'b1101100000100,
13'b1101100010100,
13'b1101100100011,
13'b1101100100100,
13'b1101100110011: edge_mask_reg_512p3[306] <= 1'b1;
 		default: edge_mask_reg_512p3[306] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b101101010,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11001001001,
13'b11001001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100001001001,
13'b100001001010,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b101001101001,
13'b101001101010,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b1000001110101,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1001001110100,
13'b1001001110101,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1011010100101,
13'b1011010100110,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100011,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110011,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100100100,
13'b1100011100011,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011110011,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010100,
13'b1100100010101,
13'b1100100010110,
13'b1100100100100,
13'b1100100100101,
13'b1101100000100,
13'b1101100010100: edge_mask_reg_512p3[307] <= 1'b1;
 		default: edge_mask_reg_512p3[307] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000101,
13'b11011000110,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100011000101,
13'b100011000110,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101011000101,
13'b101011000110,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100101,
13'b110010100110,
13'b110010110101,
13'b110010110110,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001010000001,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1010000000100,
13'b1010000000101,
13'b1010000000110,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010010001,
13'b1010010010010,
13'b1010010010011,
13'b1011000000011,
13'b1011000000100,
13'b1011000000101,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001110001,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011010000001,
13'b1011010000010,
13'b1011010000011,
13'b1011010010001,
13'b1011010010010,
13'b1011010010011,
13'b1100000000011,
13'b1100000000100,
13'b1100000000101,
13'b1100000010011,
13'b1100000010100,
13'b1100000010101,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000110010,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100001000001,
13'b1100001000010,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1100001010100,
13'b1100001100001,
13'b1100001100010,
13'b1100001100011,
13'b1100001100100,
13'b1100001110000,
13'b1100001110001,
13'b1100001110010,
13'b1100001110011,
13'b1100010000000,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010010001,
13'b1100010010010,
13'b1101000000011,
13'b1101000000100,
13'b1101000000101,
13'b1101000010011,
13'b1101000010100,
13'b1101000010101,
13'b1101000100010,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000110010,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101001000001,
13'b1101001000010,
13'b1101001000011,
13'b1101001000100,
13'b1101001010001,
13'b1101001010010,
13'b1101001010011,
13'b1101001010100,
13'b1101001100000,
13'b1101001100001,
13'b1101001100010,
13'b1101001100011,
13'b1101001110000,
13'b1101001110001,
13'b1101001110010,
13'b1101001110011,
13'b1101010000000,
13'b1101010000001,
13'b1101010000010,
13'b1101010000011,
13'b1110000000011,
13'b1110000000100,
13'b1110000000101,
13'b1110000010011,
13'b1110000010100,
13'b1110000010101,
13'b1110000100010,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000110010,
13'b1110000110011,
13'b1110000110100,
13'b1110001000001,
13'b1110001000010,
13'b1110001000011,
13'b1110001000100,
13'b1110001010001,
13'b1110001010010,
13'b1110001010011,
13'b1110001100000,
13'b1110001100001,
13'b1110001100010,
13'b1110001100011,
13'b1110001110000,
13'b1110001110001,
13'b1110001110010,
13'b1110010000000,
13'b1110010000001,
13'b1110010000010,
13'b1111000000011,
13'b1111000000100,
13'b1111000010011,
13'b1111000010100,
13'b1111000010101,
13'b1111000100010,
13'b1111000100011,
13'b1111000100100,
13'b1111000110001,
13'b1111000110010,
13'b1111000110011,
13'b1111000110100,
13'b1111001000001,
13'b1111001000010,
13'b1111001000011,
13'b1111001010000,
13'b1111001010001,
13'b1111001010010,
13'b1111001010011,
13'b1111001100000,
13'b1111001100001,
13'b1111001100010,
13'b1111001100011,
13'b1111001110000,
13'b1111001110001,
13'b1111001110010,
13'b1111010000000,
13'b1111010000001,
13'b1111010000010: edge_mask_reg_512p3[308] <= 1'b1;
 		default: edge_mask_reg_512p3[308] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011001001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111001,
13'b11010111010,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001001011,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101001,
13'b101010101010,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000011001,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1010000000011,
13'b1010000000100,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1011000110101,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100101,
13'b1011001100110: edge_mask_reg_512p3[309] <= 1'b1;
 		default: edge_mask_reg_512p3[309] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001011000,
13'b11001011001,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001001000,
13'b100001001001,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001001000,
13'b101001001001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000101000,
13'b110000101001,
13'b110000111000,
13'b110000111001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100: edge_mask_reg_512p3[310] <= 1'b1;
 		default: edge_mask_reg_512p3[310] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100001000,
13'b10100001001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b110000111000,
13'b110000111001,
13'b110001001000,
13'b110001001001,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b111001001000,
13'b111001001001,
13'b111001011000,
13'b111001011001,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001111000,
13'b111001111001,
13'b111001111010,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010101011,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111010111011,
13'b111011001001,
13'b111011001010,
13'b111011001011,
13'b1000001010111,
13'b1000001011000,
13'b1000001011001,
13'b1000001100111,
13'b1000001101000,
13'b1000001101001,
13'b1000001111000,
13'b1000001111001,
13'b1000001111010,
13'b1000010001000,
13'b1000010001001,
13'b1000010001010,
13'b1000010011000,
13'b1000010011001,
13'b1000010011010,
13'b1000010101000,
13'b1000010101001,
13'b1000010101010,
13'b1000010101011,
13'b1000010111001,
13'b1000010111010,
13'b1000010111011,
13'b1000011001001,
13'b1000011001010,
13'b1000011001011,
13'b1001001010111,
13'b1001001011000,
13'b1001001011001,
13'b1001001100111,
13'b1001001101000,
13'b1001001101001,
13'b1001001111000,
13'b1001001111001,
13'b1001001111010,
13'b1001010001000,
13'b1001010001001,
13'b1001010001010,
13'b1001010011000,
13'b1001010011001,
13'b1001010011010,
13'b1001010101000,
13'b1001010101001,
13'b1001010101010,
13'b1001010101011,
13'b1001010111001,
13'b1001010111010,
13'b1001010111011,
13'b1001011001001,
13'b1001011001010,
13'b1001011001011,
13'b1001011011010,
13'b1010001001000,
13'b1010001010111,
13'b1010001011000,
13'b1010001011001,
13'b1010001100111,
13'b1010001101000,
13'b1010001101001,
13'b1010001110111,
13'b1010001111000,
13'b1010001111001,
13'b1010001111010,
13'b1010010001000,
13'b1010010001001,
13'b1010010001010,
13'b1010010011000,
13'b1010010011001,
13'b1010010011010,
13'b1010010011011,
13'b1010010101000,
13'b1010010101001,
13'b1010010101010,
13'b1010010101011,
13'b1010010111001,
13'b1010010111010,
13'b1010010111011,
13'b1010011001001,
13'b1010011001010,
13'b1010011001011,
13'b1010011011010,
13'b1011001000111,
13'b1011001001000,
13'b1011001010111,
13'b1011001011000,
13'b1011001011001,
13'b1011001100111,
13'b1011001101000,
13'b1011001101001,
13'b1011001111000,
13'b1011001111001,
13'b1011001111010,
13'b1011010001000,
13'b1011010001001,
13'b1011010001010,
13'b1011010011000,
13'b1011010011001,
13'b1011010011010,
13'b1011010011011,
13'b1011010101001,
13'b1011010101010,
13'b1011010101011,
13'b1011010111001,
13'b1011010111010,
13'b1011010111011,
13'b1011010111100,
13'b1011011001010,
13'b1011011001011,
13'b1011011001100,
13'b1100001010111,
13'b1100001011000,
13'b1100001011001,
13'b1100001100111,
13'b1100001101000,
13'b1100001101001,
13'b1100001110111,
13'b1100001111000,
13'b1100001111001,
13'b1100001111010,
13'b1100010001000,
13'b1100010001001,
13'b1100010001010,
13'b1100010001011,
13'b1100010011000,
13'b1100010011001,
13'b1100010011010,
13'b1100010011011,
13'b1100010101001,
13'b1100010101010,
13'b1100010101011,
13'b1100010101100,
13'b1100010111001,
13'b1100010111010,
13'b1100010111011,
13'b1100010111100,
13'b1100011001010,
13'b1100011001011,
13'b1100011001100,
13'b1100011011011,
13'b1101001010111,
13'b1101001011000,
13'b1101001011001,
13'b1101001100111,
13'b1101001101000,
13'b1101001101001,
13'b1101001110111,
13'b1101001111000,
13'b1101001111001,
13'b1101001111010,
13'b1101010001000,
13'b1101010001001,
13'b1101010001010,
13'b1101010001011,
13'b1101010011000,
13'b1101010011001,
13'b1101010011010,
13'b1101010011011,
13'b1101010101001,
13'b1101010101010,
13'b1101010101011,
13'b1101010101100,
13'b1101010111001,
13'b1101010111010,
13'b1101010111011,
13'b1101010111100,
13'b1101011001010,
13'b1101011001011,
13'b1101011001100,
13'b1101011011011,
13'b1110001010111,
13'b1110001011000,
13'b1110001011001,
13'b1110001100111,
13'b1110001101000,
13'b1110001101001,
13'b1110001110110,
13'b1110001110111,
13'b1110001111000,
13'b1110001111001,
13'b1110001111010,
13'b1110010000111,
13'b1110010001000,
13'b1110010001001,
13'b1110010001010,
13'b1110010001011,
13'b1110010011000,
13'b1110010011001,
13'b1110010011010,
13'b1110010011011,
13'b1110010101001,
13'b1110010101010,
13'b1110010101011,
13'b1110010111001,
13'b1110010111010,
13'b1110010111011,
13'b1110010111100,
13'b1110011001010,
13'b1110011001011,
13'b1110011001100,
13'b1111001010111,
13'b1111001011000,
13'b1111001011001,
13'b1111001100110,
13'b1111001100111,
13'b1111001101000,
13'b1111001101001,
13'b1111001110110,
13'b1111001110111,
13'b1111001111000,
13'b1111001111001,
13'b1111001111010,
13'b1111010000111,
13'b1111010001000,
13'b1111010001001,
13'b1111010001010,
13'b1111010010111,
13'b1111010011000,
13'b1111010011001,
13'b1111010011010,
13'b1111010101000,
13'b1111010101001,
13'b1111010101010,
13'b1111010101011,
13'b1111010111001,
13'b1111010111010,
13'b1111010111011,
13'b1111011001010,
13'b1111011001011: edge_mask_reg_512p3[311] <= 1'b1;
 		default: edge_mask_reg_512p3[311] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100101000,
13'b101100101001,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001101000101,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1100101010100,
13'b1100101010101,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110001,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100110000001,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110010001,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110100001,
13'b1100110100010,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110110001,
13'b1100110110010,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111100011,
13'b1100111100100,
13'b1101101100010,
13'b1101101110010,
13'b1101101110011,
13'b1101110000010,
13'b1101110000011,
13'b1101110010001,
13'b1101110010010,
13'b1101110010011,
13'b1101110100001,
13'b1101110100010,
13'b1101110100011,
13'b1101110110001,
13'b1101110110010,
13'b1101111000001,
13'b1101111000010,
13'b1101111010001: edge_mask_reg_512p3[312] <= 1'b1;
 		default: edge_mask_reg_512p3[312] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100011,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1010110100100,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111100000,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1011110100100,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111010000,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100000,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1100110110011,
13'b1100110110100,
13'b1100111000000,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111010000,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111100011,
13'b1100111100100: edge_mask_reg_512p3[313] <= 1'b1;
 		default: edge_mask_reg_512p3[313] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101110000111,
13'b101110001000,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001110100100,
13'b1001110100101,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1010110100100,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111010000,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111100000,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111110000,
13'b1010111110001,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1011110100100,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011111000000,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111010000,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111100000,
13'b1011111100001,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1100110110011,
13'b1100110110100,
13'b1100111000001,
13'b1100111000010,
13'b1100111000011,
13'b1100111000100,
13'b1100111010000,
13'b1100111010001,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111100000,
13'b1100111100001,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111110011: edge_mask_reg_512p3[314] <= 1'b1;
 		default: edge_mask_reg_512p3[314] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011010,
13'b1100011011,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011010,
13'b10100011011,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001010,
13'b11100001011,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101010,
13'b100011101011,
13'b100011111010,
13'b100011111011,
13'b101000111001,
13'b101000111010,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b110001001000,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011011000,
13'b110011011001,
13'b111001001000,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b1000001000111,
13'b1000001001000,
13'b1000001010111,
13'b1000001011000,
13'b1000001011001,
13'b1000001100111,
13'b1000001101000,
13'b1000001101001,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000001111001,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010001001,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010111,
13'b1000011011000,
13'b1001001001000,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1001001011001,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001101001,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001001111001,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010001001,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010111,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1010001100110,
13'b1010001100111,
13'b1010001101000,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010111,
13'b1011001010110,
13'b1011001010111,
13'b1011001011000,
13'b1011001100110,
13'b1011001100111,
13'b1011001101000,
13'b1011001110110,
13'b1011001110111,
13'b1011001111000,
13'b1011010000110,
13'b1011010000111,
13'b1011010001000,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1100001010110,
13'b1100001010111,
13'b1100001011000,
13'b1100001100110,
13'b1100001100111,
13'b1100001101000,
13'b1100001110110,
13'b1100001110111,
13'b1100001111000,
13'b1100010000110,
13'b1100010000111,
13'b1100010001000,
13'b1100010010110,
13'b1100010010111,
13'b1100010011000,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1101001100111,
13'b1101001101000,
13'b1101001110110,
13'b1101001110111,
13'b1101001111000,
13'b1101010000110,
13'b1101010000111,
13'b1101010001000,
13'b1101010010110,
13'b1101010010111,
13'b1101010011000,
13'b1101010100110,
13'b1101010100111,
13'b1101010101000,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1110001100111,
13'b1110001101000,
13'b1110001110111,
13'b1110001111000,
13'b1110001111001,
13'b1110010000111,
13'b1110010001000,
13'b1110010010110,
13'b1110010010111,
13'b1110010011000,
13'b1110010100110,
13'b1110010100111,
13'b1110010101000,
13'b1110010110110,
13'b1110010110111,
13'b1110010111000,
13'b1110011000110,
13'b1110011000111,
13'b1110011001000,
13'b1111001100111,
13'b1111001101000,
13'b1111001110111,
13'b1111001111000,
13'b1111010000111,
13'b1111010001000,
13'b1111010010111: edge_mask_reg_512p3[315] <= 1'b1;
 		default: edge_mask_reg_512p3[315] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100000111,
13'b100100001000,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100000111,
13'b101100001000,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110100010111,
13'b110100011000,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010101,
13'b1000111010110,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010101,
13'b1001111010110,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1011100110011,
13'b1011100110100,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111010100,
13'b1100100110011,
13'b1100100110100,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110110100,
13'b1100110110101,
13'b1100111000100,
13'b1100111000101,
13'b1100111010100,
13'b1101101000010,
13'b1101101000011,
13'b1101101000100,
13'b1101101010010,
13'b1101101010011,
13'b1101101010100,
13'b1101101100010,
13'b1101101100011,
13'b1101101100100,
13'b1101101110011,
13'b1101101110100,
13'b1101110000011,
13'b1101110000100,
13'b1101110000101,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1101110100011,
13'b1101110100100,
13'b1101110100101,
13'b1101110110100,
13'b1101110110101,
13'b1110101000010,
13'b1110101000011,
13'b1110101000100,
13'b1110101010010,
13'b1110101010011,
13'b1110101010100,
13'b1110101100010,
13'b1110101100011,
13'b1110101100100,
13'b1110101110010,
13'b1110101110011,
13'b1110101110100,
13'b1110110000011,
13'b1110110000100,
13'b1110110000101,
13'b1110110010011,
13'b1110110010100,
13'b1110110010101,
13'b1110110100011,
13'b1110110100100,
13'b1110110100101,
13'b1110110110100,
13'b1110110110101,
13'b1111101000010,
13'b1111101000011,
13'b1111101000100,
13'b1111101010010,
13'b1111101010011,
13'b1111101010100,
13'b1111101100010,
13'b1111101100011,
13'b1111101100100,
13'b1111101110010,
13'b1111101110011,
13'b1111101110100,
13'b1111110000011,
13'b1111110000100,
13'b1111110010011,
13'b1111110010100,
13'b1111110010101,
13'b1111110100011,
13'b1111110100100,
13'b1111110100101,
13'b1111110110100,
13'b1111110110101: edge_mask_reg_512p3[316] <= 1'b1;
 		default: edge_mask_reg_512p3[316] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b1001100100,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110100,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000100,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b11001000011,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010010101,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010010101,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001100001,
13'b110001100010,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010101,
13'b111000010110,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100101,
13'b111000100110,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110101,
13'b111000110110,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000101,
13'b111001000110,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001100000,
13'b1000001100001,
13'b1001000010000,
13'b1001000010001,
13'b1001000100000,
13'b1001000100001,
13'b1001000110000,
13'b1001000110001,
13'b1001001000000,
13'b1001001000001,
13'b1001001010000,
13'b1001001010001,
13'b1001001100000,
13'b1001001100001,
13'b1010000100000,
13'b1010000110000,
13'b1010001000000,
13'b1010001000001,
13'b1010001010000: edge_mask_reg_512p3[317] <= 1'b1;
 		default: edge_mask_reg_512p3[317] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001010100,
13'b11001010101,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b101000100001,
13'b101000100010,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000100000,
13'b111000100001,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000100000,
13'b1001000010000: edge_mask_reg_512p3[318] <= 1'b1;
 		default: edge_mask_reg_512p3[318] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b11001000000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b100000110000,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000000,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010011,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110110,
13'b100001110111,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110110,
13'b101001110111,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010110,
13'b111000010111,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100110,
13'b111000100111,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110110,
13'b111000110111,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010: edge_mask_reg_512p3[319] <= 1'b1;
 		default: edge_mask_reg_512p3[319] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100101000111,
13'b100101001000,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101101000111,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b1000101110111,
13'b1000101111000,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1001101110110,
13'b1001101110111,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1010101110110,
13'b1010101110111,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1011101110110,
13'b1011101110111,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1100101110110,
13'b1100101110111,
13'b1100110000101,
13'b1100110000110,
13'b1100110000111,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1100110100100,
13'b1100110100101,
13'b1100110100110,
13'b1100110100111,
13'b1100110101000,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000011,
13'b1100111000100,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111010110,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111100110,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1101101110110,
13'b1101101110111,
13'b1101110000101,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1101110010100,
13'b1101110010101,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1101110100111,
13'b1101110101000,
13'b1101110110011,
13'b1101110110100,
13'b1101110110101,
13'b1101110110110,
13'b1101110110111,
13'b1101111000011,
13'b1101111000100,
13'b1101111000101,
13'b1101111000110,
13'b1101111000111,
13'b1101111010010,
13'b1101111010011,
13'b1101111010100,
13'b1101111010101,
13'b1101111010110,
13'b1101111100010,
13'b1101111100011,
13'b1101111100100,
13'b1101111100101,
13'b1101111110011,
13'b1101111110100,
13'b1101111110101,
13'b1110101110110,
13'b1110101110111,
13'b1110110000101,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110010100,
13'b1110110010101,
13'b1110110010110,
13'b1110110010111,
13'b1110110011000,
13'b1110110100100,
13'b1110110100101,
13'b1110110100110,
13'b1110110100111,
13'b1110110101000,
13'b1110110110011,
13'b1110110110100,
13'b1110110110101,
13'b1110110110110,
13'b1110110110111,
13'b1110111000011,
13'b1110111000100,
13'b1110111000101,
13'b1110111000110,
13'b1110111000111,
13'b1110111010010,
13'b1110111010011,
13'b1110111010100,
13'b1110111010101,
13'b1110111010110,
13'b1110111100010,
13'b1110111100011,
13'b1110111100100,
13'b1110111100101,
13'b1110111110010,
13'b1110111110011,
13'b1110111110100,
13'b1110111110101,
13'b1111101110110,
13'b1111101110111,
13'b1111110000101,
13'b1111110000110,
13'b1111110000111,
13'b1111110001000,
13'b1111110010101,
13'b1111110010110,
13'b1111110010111,
13'b1111110011000,
13'b1111110100100,
13'b1111110100101,
13'b1111110100110,
13'b1111110100111,
13'b1111110101000,
13'b1111110110011,
13'b1111110110100,
13'b1111110110101,
13'b1111110110110,
13'b1111110110111,
13'b1111111000011,
13'b1111111000100,
13'b1111111000101,
13'b1111111000110,
13'b1111111000111,
13'b1111111010010,
13'b1111111010011,
13'b1111111010100,
13'b1111111010101,
13'b1111111010110,
13'b1111111100001,
13'b1111111100010,
13'b1111111100011,
13'b1111111100100,
13'b1111111100101,
13'b1111111110010,
13'b1111111110011,
13'b1111111110100: edge_mask_reg_512p3[320] <= 1'b1;
 		default: edge_mask_reg_512p3[320] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[321] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001001100,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100000111100,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000101011,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101000111011,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001001011,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101001,
13'b101001101010,
13'b101001111001,
13'b101001111010,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001011001,
13'b111000011000,
13'b111000011001,
13'b111000011010,
13'b111000101000,
13'b111000101001,
13'b111000101010,
13'b111000111000,
13'b111000111001,
13'b111000111010,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b1000000011000,
13'b1000000011001,
13'b1000000011010,
13'b1000000100111,
13'b1000000101000,
13'b1000000101001,
13'b1000000101010,
13'b1000000110111,
13'b1000000111000,
13'b1000000111001,
13'b1000000111010,
13'b1000001000111,
13'b1000001001000,
13'b1000001001001,
13'b1000001001010,
13'b1000001011000,
13'b1001000010111,
13'b1001000011000,
13'b1001000011001,
13'b1001000011010,
13'b1001000100111,
13'b1001000101000,
13'b1001000101001,
13'b1001000101010,
13'b1001000110111,
13'b1001000111000,
13'b1001000111001,
13'b1001000111010,
13'b1001001000111,
13'b1001001001000,
13'b1001001001001,
13'b1010000001000,
13'b1010000001001,
13'b1010000010111,
13'b1010000011000,
13'b1010000011001,
13'b1010000100111,
13'b1010000101000,
13'b1010000101001,
13'b1010000101010,
13'b1010000110111,
13'b1010000111000,
13'b1010000111001,
13'b1010000111010,
13'b1010001000111,
13'b1010001001000,
13'b1010001001001,
13'b1010001011000,
13'b1011000000111,
13'b1011000001000,
13'b1011000001001,
13'b1011000010111,
13'b1011000011000,
13'b1011000011001,
13'b1011000100111,
13'b1011000101000,
13'b1011000101001,
13'b1011000110111,
13'b1011000111000,
13'b1011000111001,
13'b1011001000111,
13'b1011001001000,
13'b1011001001001,
13'b1011001010111,
13'b1011001011000,
13'b1100000000111,
13'b1100000001000,
13'b1100000001001,
13'b1100000010111,
13'b1100000011000,
13'b1100000011001,
13'b1100000100111,
13'b1100000101000,
13'b1100000101001,
13'b1100000110111,
13'b1100000111000,
13'b1100000111001,
13'b1100001000111,
13'b1100001001000,
13'b1100001001001,
13'b1100001010111,
13'b1100001011000,
13'b1101000000111,
13'b1101000001000,
13'b1101000010111,
13'b1101000011000,
13'b1101000011001,
13'b1101000100110,
13'b1101000100111,
13'b1101000101000,
13'b1101000101001,
13'b1101000110110,
13'b1101000110111,
13'b1101000111000,
13'b1101000111001,
13'b1101001000111,
13'b1101001001000,
13'b1110000000111,
13'b1110000010111,
13'b1110000011000,
13'b1110000100110,
13'b1110000100111,
13'b1110000101000,
13'b1110000110110,
13'b1110000110111,
13'b1110000111000,
13'b1110001000111,
13'b1110001001000,
13'b1111000010111,
13'b1111000011000,
13'b1111000100110,
13'b1111000100111,
13'b1111000101000,
13'b1111000110110,
13'b1111000110111,
13'b1111000111000,
13'b1111001000111: edge_mask_reg_512p3[322] <= 1'b1;
 		default: edge_mask_reg_512p3[322] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010000,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100000,
13'b11100001,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110000,
13'b11110001,
13'b11110010,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000000,
13'b100000001,
13'b100000010,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010000,
13'b100010001,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100000,
13'b100100001,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110000,
13'b100110001,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000000,
13'b101000001,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010000,
13'b101010001,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010000,
13'b1011010001,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100000,
13'b1011100001,
13'b1011100010,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110000,
13'b1011110001,
13'b1011110010,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000000,
13'b1100000001,
13'b1100000010,
13'b1100000011,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010000,
13'b1100010001,
13'b1100010010,
13'b1100010011,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100000,
13'b1100100001,
13'b1100100010,
13'b1100100011,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110000,
13'b1100110001,
13'b1100110010,
13'b1100110011,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000000,
13'b1101000001,
13'b1101000010,
13'b1101000011,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010000,
13'b1101010001,
13'b1101010010,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100000,
13'b1101100001,
13'b1101100010,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110000,
13'b1101110001,
13'b1101110010,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000000,
13'b1110000001,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011010001,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011100000,
13'b10011100001,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110000,
13'b10011110001,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000000,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010000,
13'b10100010001,
13'b10100010010,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100000,
13'b10100100001,
13'b10100100010,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110000,
13'b10100110001,
13'b10100110010,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000000,
13'b10101000001,
13'b10101000010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010000,
13'b10101010001,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100000,
13'b10101100001,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110000,
13'b10101110001,
13'b10101110010,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000000,
13'b10110000001,
13'b10110000010,
13'b10110000011,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010000,
13'b10110010001,
13'b10110010010,
13'b10110010011,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100000,
13'b10110100001,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011110000,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000000,
13'b11100000001,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010000,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100000,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110000,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000000,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010000,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000000,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100000,
13'b11110100001,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110101,
13'b11110110110,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b101011010101,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100110,
13'b110110100111,
13'b111100010101,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101010101,
13'b111101010110,
13'b111101100101,
13'b111101100110,
13'b111101110101,
13'b111101110110: edge_mask_reg_512p3[323] <= 1'b1;
 		default: edge_mask_reg_512p3[323] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010000,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100000,
13'b11100001,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110000,
13'b11110001,
13'b11110010,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000000,
13'b100000001,
13'b100000010,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010000,
13'b100010001,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100000,
13'b100100001,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110000,
13'b100110001,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000000,
13'b101000001,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010000,
13'b101010001,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010000,
13'b1011010001,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100000,
13'b1011100001,
13'b1011100010,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110000,
13'b1011110001,
13'b1011110010,
13'b1011110011,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000000,
13'b1100000001,
13'b1100000010,
13'b1100000011,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010000,
13'b1100010001,
13'b1100010010,
13'b1100010011,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100000,
13'b1100100001,
13'b1100100010,
13'b1100100011,
13'b1100100101,
13'b1100110000,
13'b1100110001,
13'b1100110010,
13'b1100110011,
13'b1100110101,
13'b1101000000,
13'b1101000001,
13'b1101000010,
13'b1101000011,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010000,
13'b1101010001,
13'b1101010010,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100000,
13'b1101100001,
13'b1101100010,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110000,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b10011010001,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100000,
13'b10011100001,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110000,
13'b10011110001,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000000,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010000,
13'b10100010001,
13'b10100010010,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100000,
13'b10100100001,
13'b10100100010,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110000,
13'b10100110001,
13'b10100110010,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000000,
13'b10101000001,
13'b10101000010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010000,
13'b10101010001,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100000,
13'b10101100001,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110000,
13'b10101110001,
13'b10101110010,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110000,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000000,
13'b11100000001,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010000,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100000,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110000,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000000,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010000,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110000,
13'b11101110001,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100000,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b101011010101,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b111100010101,
13'b111100010110,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111101000101,
13'b111101000110: edge_mask_reg_512p3[324] <= 1'b1;
 		default: edge_mask_reg_512p3[324] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111001000,
13'b101111010111,
13'b101111011000,
13'b101111011001: edge_mask_reg_512p3[325] <= 1'b1;
 		default: edge_mask_reg_512p3[325] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011010,
13'b11001001001,
13'b11001001010,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b100001001001,
13'b100001001010,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b101001101001,
13'b101001101010,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100011000,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010111,
13'b111100011000,
13'b1000001110101,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010111,
13'b1000100011000,
13'b1001001110100,
13'b1001001110101,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010111,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1011010100101,
13'b1011010100110,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100011,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110011,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1100011010011,
13'b1100011010100,
13'b1100011100011,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010100,
13'b1101011110100,
13'b1101100000100,
13'b1101100000101: edge_mask_reg_512p3[326] <= 1'b1;
 		default: edge_mask_reg_512p3[326] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b101101010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11010011001,
13'b11010011010,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100010101001,
13'b100010101010,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b101010111001,
13'b101010111010,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1011011010110,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110011,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100100100,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100010100,
13'b1100100010101,
13'b1100100010110,
13'b1100100100100,
13'b1100100100101,
13'b1101100000100,
13'b1101100000101,
13'b1101100010100: edge_mask_reg_512p3[327] <= 1'b1;
 		default: edge_mask_reg_512p3[327] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001111000,
13'b11001111001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001111000,
13'b100001111001,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001111000,
13'b101001111001,
13'b110000100001,
13'b110000100010,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000011001,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111001,
13'b111001000001,
13'b111001000010,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010010,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1011000000011,
13'b1011000000100,
13'b1011000010011,
13'b1011000010100,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1100000110100,
13'b1100001000100: edge_mask_reg_512p3[328] <= 1'b1;
 		default: edge_mask_reg_512p3[328] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001111000,
13'b101001111001,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111001,
13'b111001000001,
13'b111001000010,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010010,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000010111,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1011000000100,
13'b1011000000101,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000010110,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1100000010100,
13'b1100000010101,
13'b1100000100100,
13'b1100000100101,
13'b1100000110100,
13'b1100000110101,
13'b1100001000100: edge_mask_reg_512p3[329] <= 1'b1;
 		default: edge_mask_reg_512p3[329] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010101000,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000001,
13'b111001000010,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010010,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1010000000011,
13'b1010000000100,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1011000010011,
13'b1011000010100,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100001000010,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001010010,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1101000110100,
13'b1101000110101,
13'b1101001000100,
13'b1101001000101,
13'b1101001010100,
13'b1101001010101,
13'b1101001100100,
13'b1101001100101: edge_mask_reg_512p3[330] <= 1'b1;
 		default: edge_mask_reg_512p3[330] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001111000,
13'b11001111001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001111000,
13'b101001111001,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b111000010001,
13'b111000010010,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000011001,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000001,
13'b111001000010,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010010,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1100000000010,
13'b1100000000011,
13'b1100000000100,
13'b1100000010010,
13'b1100000010011,
13'b1100000010100,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000110011,
13'b1100000110100,
13'b1100001000100: edge_mask_reg_512p3[331] <= 1'b1;
 		default: edge_mask_reg_512p3[331] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100001,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110001,
13'b101001110010,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000001,
13'b101010000010,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010001,
13'b101010010010,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100001,
13'b110010100100,
13'b110010100101,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101001,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111001,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010100001,
13'b111010100010,
13'b111010100100,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100011,
13'b1010000000011,
13'b1010000000100,
13'b1010000010011,
13'b1010000010100,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010010011,
13'b1010010010100,
13'b1011000010011,
13'b1011000010100,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001010011,
13'b1011001010100,
13'b1011001100011,
13'b1011001100100,
13'b1011001110011,
13'b1011001110100,
13'b1100000110100,
13'b1100001000100: edge_mask_reg_512p3[332] <= 1'b1;
 		default: edge_mask_reg_512p3[332] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010111,
13'b11011000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100000,
13'b11001100001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110000,
13'b11001110001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000000,
13'b11010000001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010000,
13'b100001010001,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100000,
13'b100001100001,
13'b100001100010,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110000,
13'b100001110001,
13'b100001110010,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000000,
13'b100010000001,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010000,
13'b100010010001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000001,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010000,
13'b101010010001,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110111,
13'b101010111000,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100111,
13'b110010101000,
13'b110010110111,
13'b110010111000,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000111,
13'b111010001000,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010001,
13'b1000010010010,
13'b1000010010011,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001010000010,
13'b1001010000011,
13'b1001010010010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010011,
13'b1010000010100,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001110010,
13'b1010001110011,
13'b1011000010011,
13'b1011000010100,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001010011,
13'b1011001010100,
13'b1100000110100,
13'b1100001000100: edge_mask_reg_512p3[333] <= 1'b1;
 		default: edge_mask_reg_512p3[333] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b11001000000,
13'b11001000001,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010000,
13'b11001010001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100000,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b100000110000,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000000,
13'b100001000001,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010000,
13'b100001010001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100000,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010000,
13'b101001010001,
13'b101001010011,
13'b101001010100,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100000,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100000,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1010000000011,
13'b1010000000100,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1011000010011,
13'b1011000010100,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1100000110100,
13'b1100001000100: edge_mask_reg_512p3[334] <= 1'b1;
 		default: edge_mask_reg_512p3[334] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[335] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100011001,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b110100101001,
13'b110100111000,
13'b110100111001,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100101,
13'b110110101000,
13'b110110101001,
13'b110110111000,
13'b110110111001,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000001,
13'b111110000010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100101,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100100,
13'b1000110100101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1100101010010,
13'b1100101010011,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101110010,
13'b1100101110011: edge_mask_reg_512p3[336] <= 1'b1;
 		default: edge_mask_reg_512p3[336] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100111000,
13'b101100111001,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b110101001000,
13'b110101001001,
13'b110101011000,
13'b110101011001,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110111000,
13'b110110111001,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000001,
13'b111110000010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100101,
13'b111110100110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110100100,
13'b1011110100101,
13'b1100101100100,
13'b1100101100101,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100110000001,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110010010,
13'b1100110010011,
13'b1100110010100,
13'b1100110010101,
13'b1100110010110,
13'b1100110100100,
13'b1100110100101,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1101110000010,
13'b1101110000011,
13'b1101110000100,
13'b1101110000101,
13'b1101110010010,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1110110000010,
13'b1110110000011: edge_mask_reg_512p3[337] <= 1'b1;
 		default: edge_mask_reg_512p3[337] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100111000,
13'b101100111001,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010001,
13'b101111010010,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110111000,
13'b111110111001,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110110011,
13'b1010110110100,
13'b1011101110011,
13'b1011101110100,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110010011,
13'b1011110010100,
13'b1011110100011,
13'b1011110100100: edge_mask_reg_512p3[338] <= 1'b1;
 		default: edge_mask_reg_512p3[338] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101100111000,
13'b101100111001,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b101111011011,
13'b110101001000,
13'b110101001001,
13'b110101011000,
13'b110101011001,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111001,
13'b111110000001,
13'b111110000010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001001,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1011101110011,
13'b1011101110100,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1100111000100,
13'b1100111000101,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111100110,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110: edge_mask_reg_512p3[339] <= 1'b1;
 		default: edge_mask_reg_512p3[339] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100111,
13'b11101000,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111001000,
13'b101111001001,
13'b110100011000,
13'b110100011001,
13'b110100101000,
13'b110100101001,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100101,
13'b110110101000,
13'b110110101001,
13'b110110111000,
13'b110110111001,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000001,
13'b111110000010,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100101,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100100,
13'b1000110100101,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100011,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1100100110100,
13'b1100100110101,
13'b1100100110110,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101100110,
13'b1100101110001,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100110000100,
13'b1100110000101,
13'b1101100110101,
13'b1101101000010,
13'b1101101000011,
13'b1101101000100,
13'b1101101000101,
13'b1101101000110,
13'b1101101010010,
13'b1101101010011,
13'b1101101010100,
13'b1101101010101,
13'b1101101010110,
13'b1101101100010,
13'b1101101100011,
13'b1101101100100,
13'b1101101100101,
13'b1101101110010,
13'b1110101000011,
13'b1110101010010,
13'b1110101010011,
13'b1110101010100,
13'b1110101100010,
13'b1110101100011: edge_mask_reg_512p3[340] <= 1'b1;
 		default: edge_mask_reg_512p3[340] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111000111,
13'b100111001000,
13'b101111001000,
13'b101111010111,
13'b101111011000,
13'b101111011001: edge_mask_reg_512p3[341] <= 1'b1;
 		default: edge_mask_reg_512p3[341] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000110,
13'b10010000111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000110,
13'b11010000111,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000110,
13'b100010000111,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110110,
13'b110001110111,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1101000100000,
13'b1101000100001,
13'b1101000110000,
13'b1101000110001,
13'b1101001000000,
13'b1101001000001,
13'b1110000100000,
13'b1110000110000,
13'b1110000110001,
13'b1110001000000,
13'b1110001000001: edge_mask_reg_512p3[342] <= 1'b1;
 		default: edge_mask_reg_512p3[342] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100101,
13'b11001100110,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100101,
13'b100001100110,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100110,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000000,
13'b110001000001,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010101,
13'b110001010110,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100110,
13'b111000100111,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000110000,
13'b1000000110001,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000100000,
13'b1001000100001,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000010000,
13'b1011000000000,
13'b1011000000001,
13'b1100000000000: edge_mask_reg_512p3[343] <= 1'b1;
 		default: edge_mask_reg_512p3[343] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11101001010,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100101011010,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110101100,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100110111100,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111100100,
13'b111111100101,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110011001,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1000110101001,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111001000,
13'b1000111001001,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111100100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1001110101001,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001110111000,
13'b1001110111001,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111001000,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010110110111,
13'b1010110111000,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1011110000110,
13'b1011110000111,
13'b1011110010101,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011110110110,
13'b1011110110111,
13'b1011110111000,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111000111,
13'b1011111001000,
13'b1100110010101,
13'b1100110010110,
13'b1100110010111,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110100110,
13'b1100110100111,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101,
13'b1100110110110,
13'b1100110110111,
13'b1100111000011,
13'b1100111000100,
13'b1101110010101,
13'b1101110010110,
13'b1101110010111,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1101110100111,
13'b1101110110011,
13'b1101110110100,
13'b1101110110101,
13'b1101110110110,
13'b1101110110111,
13'b1101111000011,
13'b1101111000100,
13'b1110110010101,
13'b1110110010110,
13'b1110110010111,
13'b1110110100101,
13'b1110110100110,
13'b1110110100111,
13'b1110110110101,
13'b1110110110110,
13'b1111110010110,
13'b1111110010111,
13'b1111110100110,
13'b1111110100111: edge_mask_reg_512p3[344] <= 1'b1;
 		default: edge_mask_reg_512p3[344] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b1001100100,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110100,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000100,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b11001000011,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010010101,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010010101,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001100001,
13'b110001100010,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001100000,
13'b1000001100001,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001100000,
13'b1001001100001,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010001000000,
13'b1010001000001,
13'b1010001010000,
13'b1010001010001,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000100000,
13'b1011000100001: edge_mask_reg_512p3[345] <= 1'b1;
 		default: edge_mask_reg_512p3[345] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110101,
13'b101000110110,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010: edge_mask_reg_512p3[346] <= 1'b1;
 		default: edge_mask_reg_512p3[346] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011111000,
13'b1011111001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011001000,
13'b110011001001,
13'b110011011001,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110111,
13'b111010111000,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1001000110010,
13'b1001000110011,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110000,
13'b1010001110001,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110110,
13'b1010010110111,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001100000,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001110000,
13'b1011001110001,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000001,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1100001100001,
13'b1100001100010,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1100001110001,
13'b1100001110010,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010000110,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010010110,
13'b1100010010111,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010100111,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1101001110001,
13'b1101001110010,
13'b1101001110011,
13'b1101001110100,
13'b1101010000001,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1101010000110,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010010101,
13'b1101010010110,
13'b1101010010111,
13'b1101010100010,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010100110,
13'b1101010100111,
13'b1101010110100,
13'b1101010110101,
13'b1101010110110,
13'b1110001110010,
13'b1110010000010,
13'b1110010000011,
13'b1110010000100,
13'b1110010000101,
13'b1110010010010,
13'b1110010010011,
13'b1110010010100,
13'b1110010010101,
13'b1110010010110,
13'b1110010100011,
13'b1110010100100,
13'b1110010100101,
13'b1110010100110,
13'b1110010100111,
13'b1110010110011,
13'b1110010110100,
13'b1110010110110,
13'b1111010000011,
13'b1111010000100,
13'b1111010010011,
13'b1111010010100,
13'b1111010010101,
13'b1111010100011,
13'b1111010100100,
13'b1111010100101,
13'b1111010110100,
13'b1111010110101: edge_mask_reg_512p3[347] <= 1'b1;
 		default: edge_mask_reg_512p3[347] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100101000,
13'b100101001,
13'b100101010,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b10001010011,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001100011,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001110011,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b11001000011,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001001100,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010010,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b101000101001,
13'b101000101010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000111001,
13'b101000111010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001001,
13'b101001001010,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011001,
13'b101001011010,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101001,
13'b101011101010,
13'b101011110101,
13'b101011111010,
13'b110000110100,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001011001,
13'b110001011010,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001101001,
13'b110001101010,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111001,
13'b110001111010,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001001,
13'b110010001010,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011010,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011110100,
13'b110011110101,
13'b111001010010,
13'b111001010011,
13'b111001100010,
13'b111001100011,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b1000001110010,
13'b1000010000010,
13'b1000010000011,
13'b1000010010010,
13'b1000010010011,
13'b1000010100010,
13'b1000010100011,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1001010110011,
13'b1001011000011,
13'b1001011010011: edge_mask_reg_512p3[348] <= 1'b1;
 		default: edge_mask_reg_512p3[348] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100100000110,
13'b100100000111,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b101100000111,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010000,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010000,
13'b111101010001,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100000,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110000,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101100000,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101000101,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101010101,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110001,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100101110110,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1101101010011,
13'b1101101010100,
13'b1101101010101,
13'b1101101100011,
13'b1101101100100,
13'b1101101100101,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1101101110101,
13'b1101110000100,
13'b1101110000101: edge_mask_reg_512p3[349] <= 1'b1;
 		default: edge_mask_reg_512p3[349] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101010111,
13'b101011000,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10101101000,
13'b10101101001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101101111000,
13'b101101111001,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b101111011011,
13'b110110001000,
13'b110110001001,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110011000,
13'b110110011001,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111001,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111010111,
13'b111111011000,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b111111101000,
13'b1000110010011,
13'b1000110010100,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111000110,
13'b1000111000111,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111010101,
13'b1000111010110,
13'b1000111010111,
13'b1000111011000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1000111100101,
13'b1000111100110,
13'b1000111100111,
13'b1000111101000,
13'b1001110100011,
13'b1001110100100,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1001111000111,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1001111010101,
13'b1001111010110,
13'b1001111010111,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1001111100100,
13'b1001111100101,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1010111000110,
13'b1010111010001,
13'b1010111010010,
13'b1010111010011,
13'b1010111010100,
13'b1010111010101,
13'b1010111010110,
13'b1010111010111,
13'b1010111100001,
13'b1010111100010,
13'b1010111100011,
13'b1010111100100,
13'b1010111100101,
13'b1010111100110,
13'b1010111100111,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1010111110110,
13'b1010111110111,
13'b1011111000001,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1011111000101,
13'b1011111000110,
13'b1011111010001,
13'b1011111010010,
13'b1011111010011,
13'b1011111010100,
13'b1011111010101,
13'b1011111010110,
13'b1011111100010,
13'b1011111100011,
13'b1011111100100,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111110011,
13'b1011111110100,
13'b1011111110101,
13'b1011111110110,
13'b1011111110111,
13'b1100111010010,
13'b1100111010011,
13'b1100111010100,
13'b1100111010101,
13'b1100111010110,
13'b1100111100010,
13'b1100111100011,
13'b1100111100100,
13'b1100111100101,
13'b1100111100110,
13'b1100111110011,
13'b1100111110100,
13'b1100111110101,
13'b1100111110110,
13'b1101111010011,
13'b1101111010100,
13'b1101111100011,
13'b1101111100100,
13'b1101111110011,
13'b1101111110100: edge_mask_reg_512p3[350] <= 1'b1;
 		default: edge_mask_reg_512p3[350] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b100000110101,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001011000,
13'b100001011001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001011000,
13'b101001011001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000111000,
13'b110000111001,
13'b110001001000,
13'b110001001001,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000011000,
13'b111000011001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010001,
13'b1010000010010,
13'b1011000000001,
13'b1011000000010: edge_mask_reg_512p3[351] <= 1'b1;
 		default: edge_mask_reg_512p3[351] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000110111,
13'b100000111000,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110111,
13'b101000111000,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b1000000010010,
13'b1000000010011,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1011000000010,
13'b1011000000011: edge_mask_reg_512p3[352] <= 1'b1;
 		default: edge_mask_reg_512p3[352] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000110111,
13'b100000111000,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b110000100111,
13'b110000101000,
13'b1010000000010,
13'b1010000000011: edge_mask_reg_512p3[353] <= 1'b1;
 		default: edge_mask_reg_512p3[353] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b10010010111,
13'b10010011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000110,
13'b100110000111,
13'b101010100111,
13'b101010101000,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000110,
13'b101110000111,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b111011000100,
13'b111011000101,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b1000011000100,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1010011000010,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101010001,
13'b1010101010010,
13'b1011011010000,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100010000,
13'b1011100010010: edge_mask_reg_512p3[354] <= 1'b1;
 		default: edge_mask_reg_512p3[354] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010111,
13'b1110011000,
13'b10010010111,
13'b10010011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110000,
13'b100100110001,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000111,
13'b100110001000,
13'b101010100111,
13'b101010101000,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010000,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000111,
13'b101110001000,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000101,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b111011000100,
13'b111011000101,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100101000,
13'b111100101001,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100111000,
13'b111100111001,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001000,
13'b111101001001,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100010,
13'b111101100011,
13'b1000011000100,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010010,
13'b1000101010011,
13'b1000101100010,
13'b1000101100011,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100110010,
13'b1001100110011,
13'b1001101000010,
13'b1001101000011,
13'b1010011000010,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100010010,
13'b1010100010011,
13'b1011011010000,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011: edge_mask_reg_512p3[355] <= 1'b1;
 		default: edge_mask_reg_512p3[355] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000111,
13'b1101001000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010001,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100000,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110000,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010000,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100000,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110000,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000000,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110111,
13'b100100111000,
13'b101001100110,
13'b101001100111,
13'b101001110001,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000000,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110111,
13'b101100111000,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010000,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b111010000001,
13'b111010000010,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010110,
13'b111010010111,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000000,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010000,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b1000010010001,
13'b1000010010010,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010110000,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000011000000,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011010000,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010011,
13'b1001010100010,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100010010,
13'b1001100010011,
13'b1010011000010,
13'b1010011000011,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000010,
13'b1010100000011,
13'b1011011010000,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011110011: edge_mask_reg_512p3[356] <= 1'b1;
 		default: edge_mask_reg_512p3[356] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10101111001,
13'b10101111010,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11101111010,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100110001001,
13'b100110001010,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101110011001,
13'b101110011010,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b101111011011,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b110111011010,
13'b111110111000,
13'b111110111001,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b1000110110111,
13'b1000110111000,
13'b1000111000111,
13'b1000111001000,
13'b1000111001001,
13'b1000111010111,
13'b1000111011000,
13'b1000111011001,
13'b1000111100111,
13'b1000111101000,
13'b1000111101001,
13'b1001110110111,
13'b1001110111000,
13'b1001110111001,
13'b1001111000111,
13'b1001111001000,
13'b1001111001001,
13'b1001111010110,
13'b1001111010111,
13'b1001111011000,
13'b1001111011001,
13'b1001111100110,
13'b1001111100111,
13'b1001111101000,
13'b1001111101001,
13'b1010110110111,
13'b1010110111000,
13'b1010111000110,
13'b1010111000111,
13'b1010111001000,
13'b1010111001001,
13'b1010111010110,
13'b1010111010111,
13'b1010111011000,
13'b1010111011001,
13'b1010111100110,
13'b1010111100111,
13'b1010111101000,
13'b1010111110110,
13'b1010111110111,
13'b1010111111000,
13'b1011110110111,
13'b1011110111000,
13'b1011111000110,
13'b1011111000111,
13'b1011111001000,
13'b1011111010110,
13'b1011111010111,
13'b1011111011000,
13'b1011111100101,
13'b1011111100110,
13'b1011111100111,
13'b1011111101000,
13'b1011111110101,
13'b1011111110110,
13'b1011111110111,
13'b1011111111000,
13'b1100110110111,
13'b1100110111000,
13'b1100111000101,
13'b1100111000110,
13'b1100111000111,
13'b1100111001000,
13'b1100111010101,
13'b1100111010110,
13'b1100111010111,
13'b1100111011000,
13'b1100111100101,
13'b1100111100110,
13'b1100111100111,
13'b1100111101000,
13'b1100111110101,
13'b1100111110110,
13'b1100111110111,
13'b1100111111000,
13'b1101110110111,
13'b1101111000101,
13'b1101111000110,
13'b1101111000111,
13'b1101111001000,
13'b1101111010101,
13'b1101111010110,
13'b1101111010111,
13'b1101111011000,
13'b1101111100101,
13'b1101111100110,
13'b1101111100111,
13'b1101111110100,
13'b1101111110101,
13'b1101111110110,
13'b1101111110111,
13'b1110111000101,
13'b1110111000110,
13'b1110111010101,
13'b1110111010110,
13'b1110111010111,
13'b1110111100101,
13'b1110111100110,
13'b1110111110101,
13'b1110111110110,
13'b1111111000101,
13'b1111111000110,
13'b1111111010101,
13'b1111111010110,
13'b1111111100101,
13'b1111111100110,
13'b1111111110101,
13'b1111111110110: edge_mask_reg_512p3[357] <= 1'b1;
 		default: edge_mask_reg_512p3[357] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000111,
13'b11001001000,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000111,
13'b100001001000,
13'b101000100001,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b110000100000,
13'b110000100001,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110111,
13'b110000111000,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1010000000010,
13'b1010000000011: edge_mask_reg_512p3[358] <= 1'b1;
 		default: edge_mask_reg_512p3[358] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000111,
13'b11001001000,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000111,
13'b100001001000,
13'b101000100001,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b110000100001,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000111000,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1010000000010,
13'b1010000000011: edge_mask_reg_512p3[359] <= 1'b1;
 		default: edge_mask_reg_512p3[359] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000111,
13'b11001001000,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000111,
13'b100001001000,
13'b101000100001,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b110000100001,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000111000,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1010000000010,
13'b1010000000011: edge_mask_reg_512p3[360] <= 1'b1;
 		default: edge_mask_reg_512p3[360] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000110,
13'b101000111,
13'b101010110,
13'b101010111,
13'b101100110,
13'b101100111,
13'b1101000110,
13'b1101000111,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10101010110,
13'b10101010111,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11101010110,
13'b11101010111,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100101010110,
13'b100101010111,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110101100110,
13'b110101100111,
13'b110101110001,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010110,
13'b111110010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100110,
13'b111110100111,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110110,
13'b111110110111,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000110,
13'b111111000111,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010110,
13'b111111010111,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1001110010001,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1010111000001,
13'b1010111010001,
13'b1010111100001,
13'b1010111100010,
13'b1010111110000,
13'b1010111110001,
13'b1010111110010: edge_mask_reg_512p3[361] <= 1'b1;
 		default: edge_mask_reg_512p3[361] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000110,
13'b100110000111,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000110,
13'b101110000111,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b111010110101,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b1000010110100,
13'b1000010110101,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1001010110100,
13'b1001010110101,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101010001,
13'b1010101010010,
13'b1011010110001,
13'b1011010110011,
13'b1011010110100,
13'b1011011000001,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011010000,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100100000,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1100011000001,
13'b1100011000010,
13'b1100011000011,
13'b1100011000100,
13'b1100011010001,
13'b1100011010010,
13'b1100011010011,
13'b1100011010100,
13'b1100011100000,
13'b1100011100001,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011110000,
13'b1100011110001,
13'b1100011110011,
13'b1101011000001: edge_mask_reg_512p3[362] <= 1'b1;
 		default: edge_mask_reg_512p3[362] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100111,
13'b11100101000,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100111,
13'b100100101000,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100111,
13'b101100101000,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010111,
13'b110100011000,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010101000,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000000,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010100000,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110000,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000000,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010100000,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110000,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1010010100000,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010110000,
13'b1010010110001,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000000,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1011010100011,
13'b1011010110001,
13'b1011010110010,
13'b1011010110011,
13'b1011010110100,
13'b1011011000000,
13'b1011011000001,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011010000,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110011,
13'b1011011110100,
13'b1100010110001,
13'b1100010110011,
13'b1100010110100,
13'b1100011000001,
13'b1100011000010,
13'b1100011000011,
13'b1100011000100,
13'b1100011010001,
13'b1100011010010,
13'b1100011010011,
13'b1100011010100,
13'b1100011100001,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1101011000001: edge_mask_reg_512p3[363] <= 1'b1;
 		default: edge_mask_reg_512p3[363] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000001,
13'b10101000010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110001,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000001,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000001,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000001,
13'b100110000010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100111,
13'b100110101000,
13'b101010110111,
13'b101010111000,
13'b101011000011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000000,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010000,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000001,
13'b101110000010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010111,
13'b101110011000,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010111,
13'b110110011000,
13'b111011010001,
13'b111011010010,
13'b111011100000,
13'b111011100001,
13'b111011100010,
13'b111011100111,
13'b111011101000,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110111,
13'b111011111000,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000111,
13'b111100001000,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100111,
13'b111100101000,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110111,
13'b111100111000,
13'b111101000000,
13'b111101000001,
13'b111101000111,
13'b111101001000,
13'b111101010000,
13'b111101010001,
13'b111101010111,
13'b111101011000,
13'b111101100001,
13'b111101100111,
13'b111101101000,
13'b1000011100000,
13'b1000011100001,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000100000000,
13'b1000100000001,
13'b1000100010000,
13'b1000100010001,
13'b1000100100000,
13'b1000100100001,
13'b1000100110000,
13'b1000100110001,
13'b1000101000000,
13'b1000101000001,
13'b1000101010000,
13'b1000101010001,
13'b1001011100000,
13'b1001011100001,
13'b1001011110000,
13'b1001011110001,
13'b1001100000000,
13'b1001100000001,
13'b1001100010000,
13'b1001100010001,
13'b1001100100000,
13'b1001100100001,
13'b1001100110000,
13'b1010011110000,
13'b1010011110001,
13'b1010100000000,
13'b1010100000001: edge_mask_reg_512p3[364] <= 1'b1;
 		default: edge_mask_reg_512p3[364] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001111000,
13'b10001111001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001101000,
13'b101001101001,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001001000,
13'b110001001001,
13'b110001010011,
13'b110001011000,
13'b110001011001,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000011000,
13'b111000011001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000101000,
13'b111000101001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111001000011,
13'b111001000100,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000100011,
13'b1000000100100: edge_mask_reg_512p3[365] <= 1'b1;
 		default: edge_mask_reg_512p3[365] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100101100111,
13'b100101101000,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101101101000,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111110010111,
13'b111110011000,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110111,
13'b111110111000,
13'b111110111001,
13'b111111000111,
13'b111111001000,
13'b111111001001,
13'b111111010111,
13'b111111011000,
13'b111111011001,
13'b111111100111,
13'b111111101000,
13'b111111101001,
13'b111111101010,
13'b1000110010111,
13'b1000110011000,
13'b1000110100111,
13'b1000110101000,
13'b1000110110111,
13'b1000110111000,
13'b1000110111001,
13'b1000111000111,
13'b1000111001000,
13'b1000111001001,
13'b1000111010111,
13'b1000111011000,
13'b1000111011001,
13'b1000111011010,
13'b1000111101000,
13'b1000111101001,
13'b1000111101010,
13'b1001110010111,
13'b1001110011000,
13'b1001110100111,
13'b1001110101000,
13'b1001110101001,
13'b1001110110111,
13'b1001110111000,
13'b1001110111001,
13'b1001111000111,
13'b1001111001000,
13'b1001111001001,
13'b1001111010111,
13'b1001111011000,
13'b1001111011001,
13'b1001111011010,
13'b1001111100111,
13'b1001111101000,
13'b1001111101001,
13'b1001111101010,
13'b1010110010111,
13'b1010110011000,
13'b1010110100111,
13'b1010110101000,
13'b1010110101001,
13'b1010110110111,
13'b1010110111000,
13'b1010110111001,
13'b1010111000111,
13'b1010111001000,
13'b1010111001001,
13'b1010111001010,
13'b1010111010111,
13'b1010111011000,
13'b1010111011001,
13'b1010111011010,
13'b1010111100111,
13'b1010111101000,
13'b1010111101001,
13'b1010111101010,
13'b1010111111000,
13'b1010111111001,
13'b1010111111010,
13'b1011110010111,
13'b1011110011000,
13'b1011110100111,
13'b1011110101000,
13'b1011110101001,
13'b1011110110111,
13'b1011110111000,
13'b1011110111001,
13'b1011111000111,
13'b1011111001000,
13'b1011111001001,
13'b1011111001010,
13'b1011111010111,
13'b1011111011000,
13'b1011111011001,
13'b1011111011010,
13'b1011111100111,
13'b1011111101000,
13'b1011111101001,
13'b1011111101010,
13'b1011111111000,
13'b1011111111001,
13'b1011111111010,
13'b1100110010111,
13'b1100110011000,
13'b1100110100111,
13'b1100110101000,
13'b1100110101001,
13'b1100110110111,
13'b1100110111000,
13'b1100110111001,
13'b1100111000111,
13'b1100111001000,
13'b1100111001001,
13'b1100111001010,
13'b1100111010111,
13'b1100111011000,
13'b1100111011001,
13'b1100111011010,
13'b1100111101000,
13'b1100111101001,
13'b1100111101010,
13'b1100111111000,
13'b1100111111001,
13'b1100111111010,
13'b1100111111011,
13'b1101110010111,
13'b1101110011000,
13'b1101110100110,
13'b1101110100111,
13'b1101110101000,
13'b1101110101001,
13'b1101110110110,
13'b1101110110111,
13'b1101110111000,
13'b1101110111001,
13'b1101111000110,
13'b1101111000111,
13'b1101111001000,
13'b1101111001001,
13'b1101111001010,
13'b1101111010111,
13'b1101111011000,
13'b1101111011001,
13'b1101111011010,
13'b1101111101000,
13'b1101111101001,
13'b1101111101010,
13'b1101111111000,
13'b1101111111001,
13'b1101111111010,
13'b1101111111011,
13'b1110110010111,
13'b1110110011000,
13'b1110110100110,
13'b1110110100111,
13'b1110110101000,
13'b1110110101001,
13'b1110110110110,
13'b1110110110111,
13'b1110110111000,
13'b1110110111001,
13'b1110111000110,
13'b1110111000111,
13'b1110111001000,
13'b1110111001001,
13'b1110111001010,
13'b1110111010111,
13'b1110111011000,
13'b1110111011001,
13'b1110111011010,
13'b1110111101000,
13'b1110111101001,
13'b1110111101010,
13'b1110111111000,
13'b1110111111001,
13'b1110111111010,
13'b1110111111011,
13'b1111110010111,
13'b1111110011000,
13'b1111110100110,
13'b1111110100111,
13'b1111110101000,
13'b1111110110110,
13'b1111110110111,
13'b1111110111000,
13'b1111110111001,
13'b1111111000110,
13'b1111111000111,
13'b1111111001000,
13'b1111111001001,
13'b1111111010111,
13'b1111111011000,
13'b1111111011001,
13'b1111111011010,
13'b1111111100111,
13'b1111111101000,
13'b1111111101001,
13'b1111111101010,
13'b1111111111000,
13'b1111111111001,
13'b1111111111010: edge_mask_reg_512p3[366] <= 1'b1;
 		default: edge_mask_reg_512p3[366] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000111,
13'b11011001000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000111,
13'b101011001000,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110111,
13'b110010111000,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010110,
13'b111010010111,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010110,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010101,
13'b1001010010110,
13'b1010000000100,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010101,
13'b1010010010110,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010010100,
13'b1011010010101,
13'b1100000010010,
13'b1100000010011,
13'b1100000010100,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000110010,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100001000010,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001010010,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001100010,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1100001100110,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1100010010101,
13'b1101000010010,
13'b1101000010011,
13'b1101000010100,
13'b1101000100010,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000110010,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101001000010,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001010010,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001100010,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001110010,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1101010010100,
13'b1101010010101,
13'b1110000010010,
13'b1110000010011,
13'b1110000010100,
13'b1110000100010,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000110010,
13'b1110000110011,
13'b1110000110100,
13'b1110000110101,
13'b1110001000010,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1110001010010,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001110010,
13'b1110001110011,
13'b1110001110100,
13'b1110001110101,
13'b1110010000011,
13'b1110010000100,
13'b1110010000101,
13'b1111000010010,
13'b1111000010011,
13'b1111000100010,
13'b1111000100011,
13'b1111000100100,
13'b1111000110001,
13'b1111000110010,
13'b1111000110011,
13'b1111000110100,
13'b1111001000001,
13'b1111001000010,
13'b1111001000011,
13'b1111001000100,
13'b1111001010010,
13'b1111001010011,
13'b1111001010100,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001110010,
13'b1111001110011,
13'b1111001110100,
13'b1111010000010,
13'b1111010000011: edge_mask_reg_512p3[367] <= 1'b1;
 		default: edge_mask_reg_512p3[367] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1011000000001,
13'b1011000000010,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000010100,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1100001000011,
13'b1100001000100,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1101000010011,
13'b1101000010100,
13'b1101000100000,
13'b1101000100001,
13'b1101000100010,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000110000,
13'b1101000110001,
13'b1101000110010,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101001000000,
13'b1101001000001,
13'b1101001000010,
13'b1101001000011,
13'b1101001000100,
13'b1110000010001,
13'b1110000010010,
13'b1110000010011,
13'b1110000010100,
13'b1110000100000,
13'b1110000100001,
13'b1110000100010,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000110000,
13'b1110000110001,
13'b1110000110010,
13'b1110000110011,
13'b1110000110100,
13'b1110000110101,
13'b1110001000000,
13'b1110001000011,
13'b1110001000100,
13'b1111000010001,
13'b1111000010010,
13'b1111000010011,
13'b1111000100000,
13'b1111000100001,
13'b1111000100010,
13'b1111000100011,
13'b1111000100100,
13'b1111000110000,
13'b1111000110001,
13'b1111000110010,
13'b1111000110011,
13'b1111000110100: edge_mask_reg_512p3[368] <= 1'b1;
 		default: edge_mask_reg_512p3[368] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b101010111001,
13'b101010111010,
13'b101011000101,
13'b101011000110,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1001011010011,
13'b1001011010100,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1010011010011,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100100010,
13'b1010100100011,
13'b1011011100011,
13'b1011011100100,
13'b1011011110011,
13'b1011011110100,
13'b1011100000011: edge_mask_reg_512p3[369] <= 1'b1;
 		default: edge_mask_reg_512p3[369] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b101011010,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b11001011010,
13'b11001011011,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b100001101010,
13'b100001101011,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001010,
13'b101010001000,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110010001000,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b111010000111,
13'b111010001000,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100010100,
13'b111100010101,
13'b1000010001000,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010100,
13'b1000100010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000011,
13'b1010100000100,
13'b1011010010111,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100011,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011110011,
13'b1011011110100,
13'b1011011110101,
13'b1011100000011,
13'b1011100000100,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1100011110100,
13'b1100011110101,
13'b1101010100110,
13'b1101010100111,
13'b1101010101000,
13'b1101010110101,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000101,
13'b1101011000110,
13'b1101011000111,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011100101,
13'b1101011100110,
13'b1110010100110,
13'b1110010100111,
13'b1110010101000,
13'b1110010110110,
13'b1110010110111,
13'b1110010111000,
13'b1110011000110,
13'b1110011000111: edge_mask_reg_512p3[370] <= 1'b1;
 		default: edge_mask_reg_512p3[370] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10101001,
13'b10101010,
13'b10101011,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101010,
13'b1010101011,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011010,
13'b10010011011,
13'b10010101010,
13'b10010101011,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001001100,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011010,
13'b11010011011,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100000111100,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001001100,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101010,
13'b100001101011,
13'b100001111010,
13'b100001111011,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000011001,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110101,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000101,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001001010,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001011010,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000011000,
13'b1000000011001,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000101001,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000000111001,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1000001001001,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001011001,
13'b1000001101000,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000010111,
13'b1001000011000,
13'b1001000011001,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000101001,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001000111000,
13'b1001000111001,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001001000,
13'b1001001001001,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1001001011001,
13'b1010000000100,
13'b1010000000101,
13'b1010000000110,
13'b1010000000111,
13'b1010000001000,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000010111,
13'b1010000011000,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000101000,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010000111000,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001001000,
13'b1010001010101,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1011000000110,
13'b1011000000111,
13'b1011000010110,
13'b1011000010111,
13'b1011000011000,
13'b1011000100110,
13'b1011000100111,
13'b1011000101000,
13'b1011000110110,
13'b1011000110111,
13'b1011000111000,
13'b1011001000101,
13'b1011001000110,
13'b1011001000111,
13'b1011001001000,
13'b1011001010111,
13'b1011001011000: edge_mask_reg_512p3[371] <= 1'b1;
 		default: edge_mask_reg_512p3[371] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10101001,
13'b10101010,
13'b10101011,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101010,
13'b1010101011,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011010,
13'b10010011011,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001001100,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001010,
13'b11010001011,
13'b11010011011,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100000111100,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001001100,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101010,
13'b100001101011,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000011001,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000011000,
13'b1000000011001,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000101001,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1000001001001,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001011001,
13'b1001000010101,
13'b1001000010110,
13'b1001000010111,
13'b1001000011000,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110110,
13'b1001000110111,
13'b1001000111000,
13'b1001001000110,
13'b1001001000111,
13'b1001001001000,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1010000000100,
13'b1010000000101,
13'b1010000000110,
13'b1010000000111,
13'b1010000010101,
13'b1010000010110,
13'b1010000010111,
13'b1010000011000,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000101000,
13'b1010000110110,
13'b1010000110111,
13'b1010000111000,
13'b1010001000110,
13'b1010001000111,
13'b1010001001000,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1011000000100,
13'b1011000000101,
13'b1011000000110,
13'b1011000000111,
13'b1011000010100,
13'b1011000010101,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1011000111000,
13'b1011001000110,
13'b1011001000111,
13'b1100000000100,
13'b1100000000101,
13'b1100000000110,
13'b1100000010100,
13'b1100000010101,
13'b1100000010110,
13'b1100000010111,
13'b1100000100101,
13'b1100000100110,
13'b1100000100111,
13'b1100000110101,
13'b1100000110110,
13'b1100000110111,
13'b1100000111000,
13'b1100001000110,
13'b1100001000111,
13'b1101000000101,
13'b1101000000110,
13'b1101000010101,
13'b1101000010110,
13'b1101000010111,
13'b1101000100101,
13'b1101000100110,
13'b1101000100111,
13'b1101000110101,
13'b1101000110110,
13'b1101000110111,
13'b1101001000110,
13'b1101001000111: edge_mask_reg_512p3[372] <= 1'b1;
 		default: edge_mask_reg_512p3[372] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101001101,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101011101,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101101101,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1101111101,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10011001010,
13'b10011001011,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101001101,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101011101,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101101101,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10101111101,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111011,
13'b100011101010,
13'b100011101011,
13'b100011111010,
13'b100011111011,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b110100001000,
13'b110100001001,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b111100001000,
13'b111100001001,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101110111,
13'b1000101111000,
13'b1000101111001,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100010111,
13'b1001100011000,
13'b1001100011001,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110111,
13'b1001101111000,
13'b1001101111001,
13'b1001110000111,
13'b1001110001000,
13'b1001110001001,
13'b1010100000111,
13'b1010100001000,
13'b1010100010111,
13'b1010100011000,
13'b1010100011001,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100101001,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101110111,
13'b1010101111000,
13'b1010110000111,
13'b1010110001000,
13'b1011100000111,
13'b1011100001000,
13'b1011100010111,
13'b1011100011000,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1101100010110,
13'b1101100010111,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110110,
13'b1101101110111,
13'b1110100010110,
13'b1110100010111,
13'b1110100100110,
13'b1110100100111,
13'b1110100101000,
13'b1110100110110,
13'b1110100110111,
13'b1110100111000,
13'b1110101000110,
13'b1110101000111,
13'b1110101010111,
13'b1111100100111: edge_mask_reg_512p3[373] <= 1'b1;
 		default: edge_mask_reg_512p3[373] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b10001010001,
13'b10001010010,
13'b10001010011,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100001,
13'b10001100010,
13'b10001100011,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001110011,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000011,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b11001000001,
13'b11001000010,
13'b11001000011,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001010001,
13'b11001010010,
13'b11001010011,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100001,
13'b11001100010,
13'b11001100011,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110001,
13'b11001110010,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000001,
13'b11010000010,
13'b11010000011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001000001,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010001,
13'b100001010010,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100001,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b101000100100,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001001001,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011001,
13'b110001011010,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101001,
13'b110001101010,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001001,
13'b110010001010,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011001,
13'b110010011010,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101001,
13'b110010101010,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111001,
13'b110010111010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001001,
13'b110011010011,
13'b110011010100,
13'b110011011001,
13'b111001000011,
13'b111001000100,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111011000011,
13'b111011000100,
13'b111011010011,
13'b111011010100,
13'b1000001110011,
13'b1000001110100,
13'b1000010000011,
13'b1000010000100,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100011,
13'b1000010100100,
13'b1000010110011,
13'b1000010110100: edge_mask_reg_512p3[374] <= 1'b1;
 		default: edge_mask_reg_512p3[374] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000100110,
13'b101000100111,
13'b101000101000: edge_mask_reg_512p3[375] <= 1'b1;
 		default: edge_mask_reg_512p3[375] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101011,
13'b10101100,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100001101,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100011101,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100101101,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b100111101,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101001101,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101011101,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b1010111011,
13'b1010111100,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100001101,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100011101,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100101101,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1100111101,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101001101,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100011101,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100101101,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10100111101,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101001101,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b11011011010,
13'b11011011011,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001010,
13'b11110001011,
13'b100011111010,
13'b100011111011,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101010,
13'b100101101011,
13'b100101111010,
13'b100101111011,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b110100001001,
13'b110100001010,
13'b110100001011,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110100111011,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b111100001001,
13'b111100001010,
13'b111100001011,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b1000100001000,
13'b1000100001001,
13'b1000100001010,
13'b1000100001011,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100011010,
13'b1000100011011,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100101010,
13'b1000100101011,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000100111011,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101001011,
13'b1000101011000,
13'b1000101011001,
13'b1001100001001,
13'b1001100001010,
13'b1001100001011,
13'b1001100010111,
13'b1001100011000,
13'b1001100011001,
13'b1001100011010,
13'b1001100011011,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100101010,
13'b1001100101011,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001100111010,
13'b1001100111011,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101001010,
13'b1001101001011,
13'b1001101011000,
13'b1001101011001,
13'b1010100001001,
13'b1010100001010,
13'b1010100010111,
13'b1010100011000,
13'b1010100011001,
13'b1010100011010,
13'b1010100011011,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100101001,
13'b1010100101010,
13'b1010100101011,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010100111010,
13'b1010100111011,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101001010,
13'b1010101001011,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1011100001010,
13'b1011100010111,
13'b1011100011000,
13'b1011100011001,
13'b1011100011010,
13'b1011100011011,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100101001,
13'b1011100101010,
13'b1011100101011,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011100111001,
13'b1011100111010,
13'b1011100111011,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101001001,
13'b1011101001010,
13'b1011101001011,
13'b1011101010111,
13'b1011101011000,
13'b1100100011000,
13'b1100100011001,
13'b1100100100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100101001,
13'b1100100101010,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100100111001,
13'b1100100111010,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101001001,
13'b1101100011000,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100101001,
13'b1101100101010,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101100111001,
13'b1101100111010,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1110100101000,
13'b1110100101001,
13'b1110100110111,
13'b1110100111000,
13'b1110100111001: edge_mask_reg_512p3[376] <= 1'b1;
 		default: edge_mask_reg_512p3[376] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000000,
13'b11100000001,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010000,
13'b11100010001,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110000,
13'b100011110001,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000000,
13'b100100000001,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010000,
13'b100100010001,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100000,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100110,
13'b100101100111,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110000,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000000,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010000,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100000,
13'b101100100001,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110000,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b110010110111,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110000,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010110,
13'b110101010111,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100111,
13'b111011101000,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110111,
13'b111011111000,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000111,
13'b111100001000,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100111,
13'b111100101000,
13'b111100110000,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b1000011010001,
13'b1000011010010,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1001011100001,
13'b1001011100010,
13'b1001011110001,
13'b1001011110010,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110001,
13'b1001100110010,
13'b1010100000001,
13'b1010100000010,
13'b1010100010001,
13'b1010100010010,
13'b1010100100001,
13'b1010100100010: edge_mask_reg_512p3[377] <= 1'b1;
 		default: edge_mask_reg_512p3[377] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111011,
13'b1001111100,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001001100,
13'b11001011010,
13'b11001011011,
13'b100000111010,
13'b100000111011,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000100101,
13'b1000000100110,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000010111,
13'b1010000000100: edge_mask_reg_512p3[378] <= 1'b1;
 		default: edge_mask_reg_512p3[378] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101000,
13'b11101001,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111011000,
13'b101111011001,
13'b101111011010,
13'b110100101001,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101001011,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111001000,
13'b110111001001,
13'b110111001010,
13'b110111011000,
13'b110111011001,
13'b111100111001,
13'b111100111010,
13'b111100111011,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110001100,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110011100,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110101100,
13'b111110111001,
13'b111110111010,
13'b111110111011,
13'b111110111100,
13'b111111001010,
13'b111111001011,
13'b111111001100,
13'b1000100111010,
13'b1000100111011,
13'b1000101001001,
13'b1000101001010,
13'b1000101001011,
13'b1000101011001,
13'b1000101011010,
13'b1000101011011,
13'b1000101011100,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101101100,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1000101111100,
13'b1000110001010,
13'b1000110001011,
13'b1000110001100,
13'b1000110011010,
13'b1000110011011,
13'b1000110011100,
13'b1000110101010,
13'b1000110101011,
13'b1000110101100,
13'b1000110111010,
13'b1000110111011,
13'b1000110111100,
13'b1000111001010,
13'b1000111001011,
13'b1000111001100,
13'b1001100111010,
13'b1001100111011,
13'b1001101001010,
13'b1001101001011,
13'b1001101001100,
13'b1001101011010,
13'b1001101011011,
13'b1001101011100,
13'b1001101101010,
13'b1001101101011,
13'b1001101101100,
13'b1001101111010,
13'b1001101111011,
13'b1001101111100,
13'b1001110001010,
13'b1001110001011,
13'b1001110001100,
13'b1001110011010,
13'b1001110011011,
13'b1001110011100,
13'b1001110101010,
13'b1001110101011,
13'b1001110101100,
13'b1001110101101,
13'b1001110111010,
13'b1001110111011,
13'b1001110111100,
13'b1001110111101,
13'b1001111001010,
13'b1001111001011,
13'b1001111001100,
13'b1010100111010,
13'b1010100111011,
13'b1010100111100,
13'b1010101001010,
13'b1010101001011,
13'b1010101001100,
13'b1010101011010,
13'b1010101011011,
13'b1010101011100,
13'b1010101101010,
13'b1010101101011,
13'b1010101101100,
13'b1010101101101,
13'b1010101111010,
13'b1010101111011,
13'b1010101111100,
13'b1010101111101,
13'b1010110001010,
13'b1010110001011,
13'b1010110001100,
13'b1010110001101,
13'b1010110011010,
13'b1010110011011,
13'b1010110011100,
13'b1010110011101,
13'b1010110101011,
13'b1010110101100,
13'b1010110101101,
13'b1010110111011,
13'b1010110111100,
13'b1010110111101,
13'b1010111001011,
13'b1010111001100,
13'b1010111001101,
13'b1011100111011,
13'b1011100111100,
13'b1011101001010,
13'b1011101001011,
13'b1011101001100,
13'b1011101011010,
13'b1011101011011,
13'b1011101011100,
13'b1011101011101,
13'b1011101101010,
13'b1011101101011,
13'b1011101101100,
13'b1011101101101,
13'b1011101111011,
13'b1011101111100,
13'b1011101111101,
13'b1011110001011,
13'b1011110001100,
13'b1011110001101,
13'b1011110011011,
13'b1011110011100,
13'b1011110011101,
13'b1011110101011,
13'b1011110101100,
13'b1011110101101,
13'b1011110111011,
13'b1011110111100,
13'b1011110111101,
13'b1011111001011,
13'b1011111001100,
13'b1011111001101,
13'b1100100111011,
13'b1100100111100,
13'b1100101001010,
13'b1100101001011,
13'b1100101001100,
13'b1100101011011,
13'b1100101011100,
13'b1100101011101,
13'b1100101101011,
13'b1100101101100,
13'b1100101101101,
13'b1100101111011,
13'b1100101111100,
13'b1100101111101,
13'b1100110001011,
13'b1100110001100,
13'b1100110001101,
13'b1100110011011,
13'b1100110011100,
13'b1100110011101,
13'b1100110101011,
13'b1100110101100,
13'b1100110101101,
13'b1100110111011,
13'b1100110111100,
13'b1100110111101,
13'b1100111001100,
13'b1100111001101,
13'b1101100111011,
13'b1101100111100,
13'b1101101001011,
13'b1101101001100,
13'b1101101011010,
13'b1101101011011,
13'b1101101011100,
13'b1101101011101,
13'b1101101101010,
13'b1101101101011,
13'b1101101101100,
13'b1101101101101,
13'b1101101111010,
13'b1101101111011,
13'b1101101111100,
13'b1101101111101,
13'b1101110001011,
13'b1101110001100,
13'b1101110001101,
13'b1101110011011,
13'b1101110011100,
13'b1101110011101,
13'b1101110101011,
13'b1101110101100,
13'b1101110101101,
13'b1101110111011,
13'b1101110111100,
13'b1101110111101,
13'b1110101001010,
13'b1110101001011,
13'b1110101001100,
13'b1110101011010,
13'b1110101011011,
13'b1110101011100,
13'b1110101101010,
13'b1110101101011,
13'b1110101101100,
13'b1110101111010,
13'b1110101111011,
13'b1110101111100,
13'b1110110001010,
13'b1110110001011,
13'b1110110001100,
13'b1110110001101,
13'b1110110011011,
13'b1110110011100,
13'b1110110011101,
13'b1110110101011,
13'b1110110101100,
13'b1110110101101,
13'b1110110111011,
13'b1110110111100,
13'b1110110111101,
13'b1111101001010,
13'b1111101001011,
13'b1111101011010,
13'b1111101011011,
13'b1111101011100,
13'b1111101101010,
13'b1111101101011,
13'b1111101101100,
13'b1111101111010,
13'b1111101111011,
13'b1111101111100,
13'b1111110001010,
13'b1111110001011,
13'b1111110001100,
13'b1111110011010,
13'b1111110011011,
13'b1111110011100,
13'b1111110011101,
13'b1111110101011,
13'b1111110101100,
13'b1111110101101,
13'b1111110111011,
13'b1111110111100,
13'b1111110111101: edge_mask_reg_512p3[379] <= 1'b1;
 		default: edge_mask_reg_512p3[379] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110101,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000110,
13'b101000100110,
13'b101000100111,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110101,
13'b110011110110,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010011,
13'b111011010100,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1001001010100,
13'b1001001010101,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010001,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110000,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000001,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010010001,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010100000,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010110000,
13'b1010010110001,
13'b1010010110010,
13'b1010010110011,
13'b1010011000000,
13'b1010011000001,
13'b1010011000010,
13'b1010011000011,
13'b1010011010001,
13'b1010011010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011010000001,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010010000,
13'b1011010010001,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010100000,
13'b1011010100001,
13'b1011010100010,
13'b1011010100011,
13'b1011010110000,
13'b1011010110001,
13'b1011010110010,
13'b1011010110011,
13'b1011011000000,
13'b1011011000001,
13'b1011011000010,
13'b1011011010001,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001100010,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1100001110010,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010010000,
13'b1100010010001,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010100000,
13'b1100010100001,
13'b1100010100010,
13'b1100010100011,
13'b1100010110000,
13'b1100010110001,
13'b1100010110010,
13'b1100011000000,
13'b1100011000001,
13'b1101001010011,
13'b1101001010100,
13'b1101001100010,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001110001,
13'b1101001110010,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101010000000,
13'b1101010000001,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010010000,
13'b1101010010001,
13'b1101010010010,
13'b1101010010011,
13'b1101010100000,
13'b1101010100001,
13'b1101010100010,
13'b1101010100011,
13'b1101010110000,
13'b1101010110001,
13'b1110001010011,
13'b1110001010100,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001110001,
13'b1110001110010,
13'b1110001110011,
13'b1110001110100,
13'b1110010000000,
13'b1110010000001,
13'b1110010000010,
13'b1110010000011,
13'b1110010010000,
13'b1110010010001,
13'b1110010010010,
13'b1110010010011,
13'b1110010100000,
13'b1110010100001,
13'b1110010100010,
13'b1110010110000,
13'b1110010110001,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001110001,
13'b1111001110010,
13'b1111001110011,
13'b1111001110100,
13'b1111010000000,
13'b1111010000001,
13'b1111010000010,
13'b1111010000011,
13'b1111010010000,
13'b1111010010001,
13'b1111010010010,
13'b1111010100000,
13'b1111010100001,
13'b1111010100010,
13'b1111010110000: edge_mask_reg_512p3[380] <= 1'b1;
 		default: edge_mask_reg_512p3[380] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110110,
13'b100010110111,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110110,
13'b101010110111,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110110,
13'b110010110111,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b1000000010011,
13'b1000000010100,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110010,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1010000010010,
13'b1010000010011,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1011000010010,
13'b1011000010011,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011010000011,
13'b1011010000100,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100000110100,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1100001000011,
13'b1100001000100,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001100001,
13'b1100001100010,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1100001110010,
13'b1100001110011,
13'b1100001110100,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1101000100000,
13'b1101000100001,
13'b1101000110000,
13'b1101000110001,
13'b1101000110010,
13'b1101000110011,
13'b1101001000000,
13'b1101001000001,
13'b1101001000010,
13'b1101001000011,
13'b1101001000100,
13'b1101001010000,
13'b1101001010001,
13'b1101001010010,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001100001,
13'b1101001100010,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001110010,
13'b1101001110011,
13'b1101001110100,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1110000110000,
13'b1110000110001,
13'b1110000110010,
13'b1110001000000,
13'b1110001000001,
13'b1110001000010,
13'b1110001010000,
13'b1110001010001,
13'b1110001010010,
13'b1110001010011,
13'b1110001010100,
13'b1110001100000,
13'b1110001100001,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001110001,
13'b1110001110010,
13'b1110001110011,
13'b1110001110100,
13'b1110010000011,
13'b1111000110001,
13'b1111001000001,
13'b1111001000010,
13'b1111001010001,
13'b1111001010010,
13'b1111001010011,
13'b1111001100001,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001110001,
13'b1111001110010,
13'b1111001110011,
13'b1111001110100,
13'b1111010000010,
13'b1111010000011: edge_mask_reg_512p3[381] <= 1'b1;
 		default: edge_mask_reg_512p3[381] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110110,
13'b100010110111,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110110,
13'b101010110111,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110110,
13'b110010110111,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000010111,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1010000000101,
13'b1010000000110,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000010111,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1011000000100,
13'b1011000000101,
13'b1011000000110,
13'b1011000010100,
13'b1011000010101,
13'b1011000010110,
13'b1011000010111,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011010000011,
13'b1011010000100,
13'b1100000000100,
13'b1100000000101,
13'b1100000000110,
13'b1100000010100,
13'b1100000010101,
13'b1100000010110,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000100110,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100000110110,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001000110,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001100010,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1100001110010,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1101000000100,
13'b1101000000101,
13'b1101000000110,
13'b1101000010100,
13'b1101000010101,
13'b1101000010110,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000100110,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101000110110,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001100010,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001110010,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1110000000100,
13'b1110000000101,
13'b1110000000110,
13'b1110000010011,
13'b1110000010100,
13'b1110000010101,
13'b1110000010110,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000100110,
13'b1110000110011,
13'b1110000110100,
13'b1110000110101,
13'b1110001000010,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1110001010010,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001110010,
13'b1110001110011,
13'b1110001110100,
13'b1110010000011,
13'b1111000010011,
13'b1111000010100,
13'b1111000010101,
13'b1111000100011,
13'b1111000100100,
13'b1111000100101,
13'b1111000110011,
13'b1111000110100,
13'b1111000110101,
13'b1111001000010,
13'b1111001000011,
13'b1111001000100,
13'b1111001010010,
13'b1111001010011,
13'b1111001010100,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001110010,
13'b1111001110011,
13'b1111001110100,
13'b1111010000010,
13'b1111010000011: edge_mask_reg_512p3[382] <= 1'b1;
 		default: edge_mask_reg_512p3[382] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100111000110,
13'b100111000111,
13'b101111000111,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b1010111110010,
13'b1010111110011,
13'b1010111110100,
13'b1010111110101,
13'b1011111110010,
13'b1011111110011,
13'b1011111110100,
13'b1100111110010,
13'b1100111110011: edge_mask_reg_512p3[383] <= 1'b1;
 		default: edge_mask_reg_512p3[383] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[384] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[385] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b1010000110,
13'b1010000111,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001110011,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001100001,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010010,
13'b100010010011,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110111,
13'b100010111000,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110111,
13'b101010111000,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000000,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010010010,
13'b111010010011,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001110000,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000010000000,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1001001000010,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001110000,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1001010000000,
13'b1001010000001,
13'b1001010000010,
13'b1010001100000,
13'b1010001100001,
13'b1010001110000,
13'b1010001110001,
13'b1010001110010,
13'b1010010000000,
13'b1010010000001,
13'b1011001110001: edge_mask_reg_512p3[386] <= 1'b1;
 		default: edge_mask_reg_512p3[386] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11100111,
13'b11101000,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101001000,
13'b1101001001,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001001,
13'b100010001001,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b110010101001,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010111000,
13'b110010111001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100011000,
13'b110100011001,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b1000010110011,
13'b1000010110100,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000001,
13'b1000100000010,
13'b1001011000001,
13'b1001011000010,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011110001,
13'b1001011110010,
13'b1010011010010,
13'b1010011100010: edge_mask_reg_512p3[387] <= 1'b1;
 		default: edge_mask_reg_512p3[387] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b11010011001,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b101010101000,
13'b101010101001,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000000,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010000,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110011000,
13'b101110011001,
13'b110010111000,
13'b110010111001,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011001000,
13'b110011001001,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100101000,
13'b110100101001,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100111000,
13'b110100111001,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101001000,
13'b110101001001,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101011000,
13'b110101011001,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101101000,
13'b110101101001,
13'b110101111000,
13'b110101111001,
13'b110110001000,
13'b110110001001,
13'b111011000011,
13'b111011000100,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100101000,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100111000,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101001000,
13'b111101001001,
13'b111101010000,
13'b111101010001,
13'b111101011000,
13'b111101011001,
13'b1000011100001,
13'b1000011100010,
13'b1000011110001,
13'b1000011110010,
13'b1000100000001,
13'b1000100010001,
13'b1000100100001: edge_mask_reg_512p3[388] <= 1'b1;
 		default: edge_mask_reg_512p3[388] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110101,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110101,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101111000,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b100010100110,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100111,
13'b100101101000,
13'b101010100110,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100111,
13'b101101101000,
13'b110010110110,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010111,
13'b110101011000,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1011011010001,
13'b1011011010010,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100100000,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1100011100010,
13'b1100011100011,
13'b1100011110000,
13'b1100011110001,
13'b1100011110010,
13'b1100011110011,
13'b1100011110100,
13'b1100100000000,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100000100,
13'b1100100010000,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100000,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1101100000000,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100000100,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100010100,
13'b1101100100001,
13'b1101100100010,
13'b1101100100011,
13'b1101100100100,
13'b1101100110011,
13'b1101100110100,
13'b1110100010001,
13'b1110100100001,
13'b1110100100010: edge_mask_reg_512p3[389] <= 1'b1;
 		default: edge_mask_reg_512p3[389] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000100,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010100,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100110,
13'b1011100111,
13'b1011110111,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b100010100110,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000001,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100000,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b101010100110,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110000,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000000,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010000,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110000,
13'b101100110001,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010101,
13'b101101010110,
13'b110010110110,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110000,
13'b110100110001,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b111011010000,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011100000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100110000,
13'b1000011010000,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100110000,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100100000,
13'b1001100100001,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1011011010001,
13'b1011011010010,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011100000001,
13'b1011100000010,
13'b1011100010001,
13'b1011100010010: edge_mask_reg_512p3[390] <= 1'b1;
 		default: edge_mask_reg_512p3[390] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110101,
13'b11101110110,
13'b100010100110,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101110101,
13'b100101110110,
13'b101010100110,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100000,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101110101,
13'b101101110110,
13'b110010110110,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100101,
13'b110101100110,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101010000,
13'b111101010001,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010101000000,
13'b1010101000001,
13'b1011011010001,
13'b1011011010010,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100010001,
13'b1011100010010: edge_mask_reg_512p3[391] <= 1'b1;
 		default: edge_mask_reg_512p3[391] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b100000110000,
13'b100000110001,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000000,
13'b100001000001,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010001,
13'b100001010010,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100001,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100101,
13'b100010100110,
13'b101000100000,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110000,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010100101,
13'b101010100110,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110000,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000000,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010101,
13'b110010010110,
13'b110010100101,
13'b110010100110,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010110,
13'b111000010111,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100110,
13'b111000100111,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110110,
13'b111000110111,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000110,
13'b111001000111,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010110,
13'b111001010111,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100110,
13'b111001100111,
13'b111001110000,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111010000000,
13'b111010000001,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001110000,
13'b1000001110001,
13'b1001000010000,
13'b1001000010001,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001110000,
13'b1010000110000,
13'b1010000110001,
13'b1010001000000,
13'b1010001000001,
13'b1010001010000,
13'b1010001010001: edge_mask_reg_512p3[392] <= 1'b1;
 		default: edge_mask_reg_512p3[392] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101100101,
13'b101100110,
13'b101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b110111010111,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b111111010110,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100011,
13'b111111100100,
13'b111111100101,
13'b111111100110,
13'b111111100111,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111010011,
13'b1000111100000,
13'b1000111100001,
13'b1000111100010,
13'b1000111100011,
13'b1000111100100,
13'b1001110100000,
13'b1001110100001,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111010000,
13'b1001111010001,
13'b1001111010010,
13'b1001111010011,
13'b1001111100000,
13'b1001111100001,
13'b1001111100010,
13'b1001111100011,
13'b1010110110000,
13'b1010110110001,
13'b1010111000000,
13'b1010111000001,
13'b1010111010000,
13'b1010111010001,
13'b1010111100000,
13'b1010111100001,
13'b1010111110000,
13'b1010111110001,
13'b1010111110010: edge_mask_reg_512p3[393] <= 1'b1;
 		default: edge_mask_reg_512p3[393] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100101000,
13'b100100101001,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010111,
13'b110111011000,
13'b111101011001,
13'b111101011010,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b1000101011001,
13'b1000101011010,
13'b1000101101000,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101110111,
13'b1000101111000,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1000110001010,
13'b1000110001011,
13'b1000110010110,
13'b1000110010111,
13'b1000110011000,
13'b1000110011001,
13'b1000110011010,
13'b1000110100110,
13'b1000110100111,
13'b1000110101000,
13'b1001101011001,
13'b1001101011010,
13'b1001101011011,
13'b1001101101000,
13'b1001101101001,
13'b1001101101010,
13'b1001101101011,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001101111001,
13'b1001101111010,
13'b1001101111011,
13'b1001101111100,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110001001,
13'b1001110001010,
13'b1001110001011,
13'b1001110001100,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1001110011001,
13'b1001110011010,
13'b1001110011011,
13'b1001110100110,
13'b1001110100111,
13'b1001110101000,
13'b1010101011001,
13'b1010101011010,
13'b1010101011011,
13'b1010101101000,
13'b1010101101001,
13'b1010101101010,
13'b1010101101011,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010101111001,
13'b1010101111010,
13'b1010101111011,
13'b1010101111100,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110001001,
13'b1010110001010,
13'b1010110001011,
13'b1010110001100,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1010110011001,
13'b1010110011010,
13'b1010110011011,
13'b1010110100110,
13'b1010110100111,
13'b1010110101000,
13'b1010110101001,
13'b1011101011010,
13'b1011101011011,
13'b1011101101000,
13'b1011101101001,
13'b1011101101010,
13'b1011101101011,
13'b1011101101100,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1011101111001,
13'b1011101111010,
13'b1011101111011,
13'b1011101111100,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1011110001001,
13'b1011110001010,
13'b1011110001011,
13'b1011110001100,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1011110011001,
13'b1011110011010,
13'b1011110011011,
13'b1011110100110,
13'b1011110100111,
13'b1011110101000,
13'b1011110101001,
13'b1100101011010,
13'b1100101011011,
13'b1100101101000,
13'b1100101101001,
13'b1100101101010,
13'b1100101101011,
13'b1100101101100,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100101111001,
13'b1100101111010,
13'b1100101111011,
13'b1100101111100,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1100110001001,
13'b1100110001010,
13'b1100110001011,
13'b1100110001100,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1100110011001,
13'b1100110011010,
13'b1100110011011,
13'b1100110100110,
13'b1100110100111,
13'b1100110101000,
13'b1100110101001,
13'b1101101011010,
13'b1101101011011,
13'b1101101101000,
13'b1101101101001,
13'b1101101101010,
13'b1101101101011,
13'b1101101101100,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101101111001,
13'b1101101111010,
13'b1101101111011,
13'b1101101111100,
13'b1101110000101,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1101110001001,
13'b1101110001010,
13'b1101110001011,
13'b1101110001100,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1101110011001,
13'b1101110011010,
13'b1101110011011,
13'b1101110100110,
13'b1101110100111,
13'b1101110101000,
13'b1101110101001,
13'b1110101011010,
13'b1110101011011,
13'b1110101101000,
13'b1110101101001,
13'b1110101101010,
13'b1110101101011,
13'b1110101101100,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110101111001,
13'b1110101111010,
13'b1110101111011,
13'b1110101111100,
13'b1110110000101,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110001001,
13'b1110110001010,
13'b1110110001011,
13'b1110110001100,
13'b1110110010110,
13'b1110110010111,
13'b1110110011000,
13'b1110110011001,
13'b1110110011010,
13'b1110110011011,
13'b1110110100110,
13'b1110110100111,
13'b1110110101000,
13'b1110110101001,
13'b1111101101000,
13'b1111101101001,
13'b1111101101010,
13'b1111101101011,
13'b1111101101100,
13'b1111101110110,
13'b1111101110111,
13'b1111101111000,
13'b1111101111001,
13'b1111101111010,
13'b1111101111011,
13'b1111101111100,
13'b1111101111101,
13'b1111110000110,
13'b1111110000111,
13'b1111110001000,
13'b1111110001001,
13'b1111110001010,
13'b1111110001011,
13'b1111110001100,
13'b1111110010110,
13'b1111110010111,
13'b1111110011000,
13'b1111110011001,
13'b1111110011010,
13'b1111110100110,
13'b1111110100111,
13'b1111110101000,
13'b1111110101001: edge_mask_reg_512p3[394] <= 1'b1;
 		default: edge_mask_reg_512p3[394] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110110,
13'b100110111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110110,
13'b1100110111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b100001000101,
13'b100001000110,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100110,
13'b100100100111,
13'b101001000101,
13'b101001000110,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100110,
13'b101100100111,
13'b110001010101,
13'b110001010110,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100110,
13'b110100100111,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b1000001110100,
13'b1000001110101,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1001001110100,
13'b1001001110101,
13'b1001010000100,
13'b1001010000101,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100101,
13'b1010011100110,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011110101,
13'b1011011110110,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010001,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010100001,
13'b1100010100010,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010110001,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100011000010,
13'b1100011000011,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011010010,
13'b1100011010011,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1100011110101,
13'b1100011110110,
13'b1101001110011,
13'b1101001110100,
13'b1101010000001,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1101010010001,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010010101,
13'b1101010100001,
13'b1101010100010,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010110001,
13'b1101010110010,
13'b1101010110011,
13'b1101010110100,
13'b1101010110101,
13'b1101010110110,
13'b1101011000010,
13'b1101011000011,
13'b1101011000100,
13'b1101011000101,
13'b1101011000110,
13'b1101011010010,
13'b1101011010011,
13'b1101011010100,
13'b1101011010101,
13'b1101011010110,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011100101,
13'b1101011100110,
13'b1101011110011,
13'b1101011110100,
13'b1101011110101,
13'b1101011110110,
13'b1110001110011,
13'b1110001110100,
13'b1110010000001,
13'b1110010000010,
13'b1110010000011,
13'b1110010000100,
13'b1110010000101,
13'b1110010010001,
13'b1110010010010,
13'b1110010010011,
13'b1110010010100,
13'b1110010010101,
13'b1110010100001,
13'b1110010100010,
13'b1110010100011,
13'b1110010100100,
13'b1110010100101,
13'b1110010110001,
13'b1110010110010,
13'b1110010110011,
13'b1110010110100,
13'b1110010110101,
13'b1110010110110,
13'b1110011000010,
13'b1110011000011,
13'b1110011000100,
13'b1110011000101,
13'b1110011000110,
13'b1110011010010,
13'b1110011010011,
13'b1110011010100,
13'b1110011010101,
13'b1110011010110,
13'b1110011100010,
13'b1110011100011,
13'b1110011100100,
13'b1110011100101,
13'b1110011100110,
13'b1110011110010,
13'b1110011110011,
13'b1110011110100,
13'b1110011110101,
13'b1110011110110,
13'b1111010000011,
13'b1111010000100,
13'b1111010010001,
13'b1111010010010,
13'b1111010010011,
13'b1111010010100,
13'b1111010010101,
13'b1111010100001,
13'b1111010100010,
13'b1111010100011,
13'b1111010100100,
13'b1111010100101,
13'b1111010110001,
13'b1111010110010,
13'b1111010110011,
13'b1111010110100,
13'b1111010110101,
13'b1111011000010,
13'b1111011000011,
13'b1111011000100,
13'b1111011000101,
13'b1111011000110,
13'b1111011010010,
13'b1111011010011,
13'b1111011010100,
13'b1111011010101,
13'b1111011010110,
13'b1111011100010,
13'b1111011100011,
13'b1111011100100,
13'b1111011100101,
13'b1111011100110,
13'b1111011110011,
13'b1111011110101,
13'b1111011110110: edge_mask_reg_512p3[395] <= 1'b1;
 		default: edge_mask_reg_512p3[395] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100011001000,
13'b100011001001,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b110011101000,
13'b110011101001,
13'b110011111000,
13'b110011111001,
13'b110100001000,
13'b110100001001,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b111011111000,
13'b111011111001,
13'b111100001000,
13'b111100001001,
13'b111100011000,
13'b111100011001,
13'b111100101000,
13'b111100101001,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b1000100001000,
13'b1000100001001,
13'b1000100001010,
13'b1000100011000,
13'b1000100011001,
13'b1000100011010,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101110111,
13'b1000101111000,
13'b1000101111001,
13'b1000110000111,
13'b1000110001000,
13'b1000110010111,
13'b1000110011000,
13'b1001011111000,
13'b1001100001000,
13'b1001100001001,
13'b1001100001010,
13'b1001100011000,
13'b1001100011001,
13'b1001100011010,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001101111001,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1010011111000,
13'b1010011111001,
13'b1010100001000,
13'b1010100001001,
13'b1010100001010,
13'b1010100011000,
13'b1010100011001,
13'b1010100011010,
13'b1010100100111,
13'b1010100101000,
13'b1010100101001,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1011011111000,
13'b1011011111001,
13'b1011100001000,
13'b1011100001001,
13'b1011100001010,
13'b1011100011000,
13'b1011100011001,
13'b1011100011010,
13'b1011100100111,
13'b1011100101000,
13'b1011100101001,
13'b1011100110111,
13'b1011100111000,
13'b1011100111001,
13'b1011101000111,
13'b1011101001000,
13'b1011101001001,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101011001,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1100011111000,
13'b1100011111001,
13'b1100100001000,
13'b1100100001001,
13'b1100100001010,
13'b1100100011000,
13'b1100100011001,
13'b1100100011010,
13'b1100100100111,
13'b1100100101000,
13'b1100100101001,
13'b1100100101010,
13'b1100100110111,
13'b1100100111000,
13'b1100100111001,
13'b1100101000111,
13'b1100101001000,
13'b1100101001001,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101011001,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101101001,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1101011111001,
13'b1101100001000,
13'b1101100001001,
13'b1101100001010,
13'b1101100011000,
13'b1101100011001,
13'b1101100011010,
13'b1101100100111,
13'b1101100101000,
13'b1101100101001,
13'b1101100101010,
13'b1101100110111,
13'b1101100111000,
13'b1101100111001,
13'b1101101000111,
13'b1101101001000,
13'b1101101001001,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101011001,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1110011111001,
13'b1110100001000,
13'b1110100001001,
13'b1110100001010,
13'b1110100011000,
13'b1110100011001,
13'b1110100011010,
13'b1110100100111,
13'b1110100101000,
13'b1110100101001,
13'b1110100101010,
13'b1110100110111,
13'b1110100111000,
13'b1110100111001,
13'b1110101000111,
13'b1110101001000,
13'b1110101001001,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101011001,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110010110,
13'b1110110010111,
13'b1110110011000,
13'b1111100001000,
13'b1111100001001,
13'b1111100001010,
13'b1111100011000,
13'b1111100011001,
13'b1111100011010,
13'b1111100100111,
13'b1111100101000,
13'b1111100101001,
13'b1111100110111,
13'b1111100111000,
13'b1111100111001,
13'b1111101000111,
13'b1111101001000,
13'b1111101001001,
13'b1111101010110,
13'b1111101010111,
13'b1111101011000,
13'b1111101011001,
13'b1111101100110,
13'b1111101100111,
13'b1111101101000,
13'b1111101110110,
13'b1111101110111,
13'b1111101111000,
13'b1111110000110,
13'b1111110000111,
13'b1111110001000,
13'b1111110010110,
13'b1111110010111: edge_mask_reg_512p3[396] <= 1'b1;
 		default: edge_mask_reg_512p3[396] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100011111000,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b111100100111,
13'b111100101000,
13'b111100110111,
13'b111100111000,
13'b111101000111,
13'b111101001000,
13'b111101010111,
13'b111101011000,
13'b111101100111,
13'b111101101000,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010111,
13'b111110011000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110111,
13'b1000101111000,
13'b1000110000111,
13'b1000110001000,
13'b1000110010111,
13'b1000110011000,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1010100100111,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1011100100110,
13'b1011100100111,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1101100100111,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1110100110101,
13'b1110100110110,
13'b1110100110111,
13'b1110101000101,
13'b1110101000110,
13'b1110101000111,
13'b1110101010101,
13'b1110101010110,
13'b1110101010111,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110010110,
13'b1110110010111,
13'b1111100110101,
13'b1111100110110,
13'b1111100110111,
13'b1111101000101,
13'b1111101000110,
13'b1111101000111,
13'b1111101010101,
13'b1111101010110,
13'b1111101010111,
13'b1111101100101,
13'b1111101100110,
13'b1111101100111,
13'b1111101110110,
13'b1111101110111,
13'b1111110000110,
13'b1111110000111,
13'b1111110010110,
13'b1111110010111: edge_mask_reg_512p3[397] <= 1'b1;
 		default: edge_mask_reg_512p3[397] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101000,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b110100101000,
13'b110100101001,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b111100111000,
13'b111100111001,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101110111,
13'b1000101111000,
13'b1000101111001,
13'b1000110000111,
13'b1000110001000,
13'b1000110010111,
13'b1000110011000,
13'b1001100111000,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001101111001,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1100100110111,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1101100110111,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1110100110111,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110010110,
13'b1110110010111,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111,
13'b1111101011000,
13'b1111101100110,
13'b1111101100111,
13'b1111101101000,
13'b1111101110110,
13'b1111101110111,
13'b1111110000110,
13'b1111110000111,
13'b1111110010110,
13'b1111110010111: edge_mask_reg_512p3[398] <= 1'b1;
 		default: edge_mask_reg_512p3[398] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100100010111,
13'b100100011000,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100010111,
13'b101100011000,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010111,
13'b111110011000,
13'b1000101000110,
13'b1000101000111,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000110,
13'b1000110000111,
13'b1000110001000,
13'b1000110010111,
13'b1000110011000,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110101,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100101,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110101,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100110000101,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1101101000101,
13'b1101101000110,
13'b1101101010100,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101100100,
13'b1101101100101,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110101,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101110000101,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1110101000101,
13'b1110101000110,
13'b1110101010100,
13'b1110101010101,
13'b1110101010110,
13'b1110101010111,
13'b1110101100100,
13'b1110101100101,
13'b1110101100110,
13'b1110101100111,
13'b1110101110100,
13'b1110101110101,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110110000101,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110010110,
13'b1110110010111,
13'b1111101010100,
13'b1111101010101,
13'b1111101010110,
13'b1111101100011,
13'b1111101100100,
13'b1111101100101,
13'b1111101100110,
13'b1111101100111,
13'b1111101110100,
13'b1111101110101,
13'b1111101110110,
13'b1111101110111,
13'b1111110000101,
13'b1111110000110,
13'b1111110000111,
13'b1111110010110,
13'b1111110010111: edge_mask_reg_512p3[399] <= 1'b1;
 		default: edge_mask_reg_512p3[399] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100001000,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b110100011000,
13'b110100011001,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b111100111000,
13'b111100111001,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101110111,
13'b1000101111000,
13'b1000101111001,
13'b1000110000111,
13'b1000110001000,
13'b1000110010111,
13'b1000110011000,
13'b1001100111000,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001101111001,
13'b1001110000110,
13'b1001110000111,
13'b1001110001000,
13'b1001110010110,
13'b1001110010111,
13'b1001110011000,
13'b1010100110111,
13'b1010100111000,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010101111001,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1010110010110,
13'b1010110010111,
13'b1010110011000,
13'b1011100110111,
13'b1011100111000,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101011001,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1011101111001,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1011110010110,
13'b1011110010111,
13'b1011110011000,
13'b1100100110111,
13'b1100100111000,
13'b1100101000111,
13'b1100101001000,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101101001,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1101100110111,
13'b1101100111000,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101011001,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101101001,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1110100110111,
13'b1110100111000,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101011001,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110010110,
13'b1110110010111,
13'b1110110011000,
13'b1111101000111,
13'b1111101001000,
13'b1111101010110,
13'b1111101010111,
13'b1111101011000,
13'b1111101100110,
13'b1111101100111,
13'b1111101101000,
13'b1111101110110,
13'b1111101110111,
13'b1111101111000,
13'b1111110000110,
13'b1111110000111,
13'b1111110001000,
13'b1111110010110,
13'b1111110010111: edge_mask_reg_512p3[400] <= 1'b1;
 		default: edge_mask_reg_512p3[400] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[401] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000110,
13'b100001000111,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000110,
13'b101001000111,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110110,
13'b110000110111,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010010,
13'b1100000010011,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011: edge_mask_reg_512p3[402] <= 1'b1;
 		default: edge_mask_reg_512p3[402] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10001010101,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010101,
13'b100001010110,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000101,
13'b101001000110,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000101,
13'b110001000110,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100011,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100011,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000100010,
13'b1001000100011,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100010,
13'b1010000100011,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000100001,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1101000010011,
13'b1110000000000,
13'b1110000000001,
13'b1110000010000: edge_mask_reg_512p3[403] <= 1'b1;
 		default: edge_mask_reg_512p3[403] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110101,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000000,
13'b1101000001,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010000,
13'b1101010001,
13'b1101010010,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100000,
13'b1101100001,
13'b1101100010,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110000,
13'b1101110001,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000000,
13'b1110000001,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110000,
13'b10100110001,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000000,
13'b10101000001,
13'b10101000010,
13'b10101000011,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010000,
13'b10101010001,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100000,
13'b10101100001,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110000,
13'b10101110001,
13'b10101110010,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000000,
13'b10110000001,
13'b10110000010,
13'b10110000011,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010000,
13'b10110010001,
13'b10110010010,
13'b10110010011,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100000,
13'b10110100001,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100000,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110000,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000000,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010000,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000000,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010000,
13'b100100010001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100000,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110000,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000101,
13'b100111000110,
13'b101011010110,
13'b101011010111,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010000,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100000,
13'b101110100001,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000101,
13'b101111000110,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110101,
13'b110110110110,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000111,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000110,
13'b111101000111,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110000,
13'b111101110001,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000101,
13'b111110000110,
13'b1000011110001,
13'b1000011110010,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101100000,
13'b1000101100001,
13'b1001100000001,
13'b1001100000010,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000001,
13'b1001101000010,
13'b1010100010000,
13'b1010100100000: edge_mask_reg_512p3[404] <= 1'b1;
 		default: edge_mask_reg_512p3[404] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010101,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110101,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000000,
13'b1101000001,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010000,
13'b1101010001,
13'b1101010010,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100000,
13'b1101100001,
13'b1101100010,
13'b1101110000,
13'b1101110001,
13'b1110000000,
13'b1110000001,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000000,
13'b10101000001,
13'b10101000010,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010000,
13'b10101010001,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100000,
13'b10101100001,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110000,
13'b10101110001,
13'b10101110010,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000000,
13'b10110000001,
13'b10110000010,
13'b10110000011,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010000,
13'b10110010001,
13'b10110010010,
13'b10110010011,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100000,
13'b10110100001,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000000,
13'b11101000001,
13'b11101000010,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010000,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000000,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110110000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b100100100110,
13'b100100100111,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110000,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101100100110,
13'b101100100111,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100000,
13'b110110100001,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b111101000001,
13'b111101000010,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b1000101010001,
13'b1000101010010,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1001101100001,
13'b1001101100010,
13'b1001101110001,
13'b1001101110010,
13'b1001110000001,
13'b1001110000010,
13'b1001110010001,
13'b1001110010010: edge_mask_reg_512p3[405] <= 1'b1;
 		default: edge_mask_reg_512p3[405] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000000,
13'b1101000001,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010000,
13'b1101010001,
13'b1101010010,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100000,
13'b1101100001,
13'b1101100010,
13'b1101110000,
13'b1101110001,
13'b1101110110,
13'b1101110111,
13'b1110000000,
13'b1110000001,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110000,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000000,
13'b10101000001,
13'b10101000010,
13'b10101000011,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010000,
13'b10101010001,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100000,
13'b10101100001,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110000,
13'b10101110001,
13'b10101110010,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000000,
13'b10110000001,
13'b10110000010,
13'b10110000011,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010000,
13'b10110010001,
13'b10110010010,
13'b10110010011,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100000,
13'b10110100001,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110000,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000000,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101010000,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000000,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100001,
13'b100100100010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110000,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000101,
13'b100111000110,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100000,
13'b101110100001,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000101,
13'b101111000110,
13'b110100010110,
13'b110100100000,
13'b110100100001,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110101,
13'b110110110110,
13'b111101000000,
13'b111101000001,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101010000,
13'b111101010001,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000000,
13'b111110000101,
13'b111110000110: edge_mask_reg_512p3[406] <= 1'b1;
 		default: edge_mask_reg_512p3[406] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000000,
13'b1101000001,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010000,
13'b1101010001,
13'b1101010010,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100000,
13'b1101100001,
13'b1101100010,
13'b1101100110,
13'b1101100111,
13'b1101110000,
13'b1101110001,
13'b1101110110,
13'b1110000000,
13'b1110000001,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000000,
13'b10101000001,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010000,
13'b10101010001,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100000,
13'b10101100001,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110000,
13'b10101110001,
13'b10101110010,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000000,
13'b10110000001,
13'b10110000010,
13'b10110000011,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010000,
13'b10110010001,
13'b10110010010,
13'b10110010011,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100000,
13'b10110100001,
13'b10110100011,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000000,
13'b11101000001,
13'b11101000010,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010000,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000000,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110000,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000000,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101010000,
13'b101101010001,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110000,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b111101100101,
13'b111101100110,
13'b111101110101,
13'b111101110110,
13'b111110000101,
13'b111110000110,
13'b111110010101,
13'b111110010110: edge_mask_reg_512p3[407] <= 1'b1;
 		default: edge_mask_reg_512p3[407] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110101,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110101,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100101,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000000,
13'b1101000001,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010000,
13'b1101010001,
13'b1101010010,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100000,
13'b1101100001,
13'b1101100010,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110000,
13'b1101110001,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000000,
13'b1110000001,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110000,
13'b10100110001,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000000,
13'b10101000001,
13'b10101000010,
13'b10101000011,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010000,
13'b10101010001,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100000,
13'b10101100001,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110000,
13'b10101110001,
13'b10101110010,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000000,
13'b10110000001,
13'b10110000010,
13'b10110000011,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110010000,
13'b10110010001,
13'b10110010010,
13'b10110010011,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100000,
13'b10110100001,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100010,
13'b11100100011,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110000,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000000,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010000,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101100000,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101110000,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000000,
13'b11110000001,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110010000,
13'b11110010001,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100000,
13'b11110100001,
13'b11110100010,
13'b11110100011,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110000,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010010,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100000,
13'b100100100001,
13'b100100100010,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110000,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000000,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010000,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100000,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100000,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110000,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000101,
13'b100111000110,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010000,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010000,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100000,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110100000,
13'b101110100001,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000101,
13'b101111000110,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110010,
13'b110011110011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110010000,
13'b110110010001,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110101,
13'b110110110110,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000111,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101100000,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101110000,
13'b111101110001,
13'b111101110010,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000101,
13'b111110000110,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101010001,
13'b1001101010010,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010101000010,
13'b1011100010000: edge_mask_reg_512p3[408] <= 1'b1;
 		default: edge_mask_reg_512p3[408] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[409] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[410] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100100,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110100,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000100,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010100,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100011,
13'b10110100100,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100011,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110001,
13'b11110110010,
13'b11110110011,
13'b11110110100,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110100001,
13'b100110100010,
13'b100110100011,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110110000,
13'b100110110001,
13'b100110110010,
13'b100110110011,
13'b100110110100,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000000,
13'b100111000001,
13'b100111000010,
13'b100111000011,
13'b100111000100,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101101010101,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000011,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010011,
13'b101111010100,
13'b101111010101,
13'b101111010110,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010110,
13'b111101110001,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000101,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010101,
13'b111111100000,
13'b111111100001,
13'b111111100010,
13'b111111100101,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111010000,
13'b1000111010001,
13'b1000111010010,
13'b1000111100000,
13'b1000111100001,
13'b1001110000000,
13'b1001110000001,
13'b1001110010000,
13'b1001110010001,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111010000,
13'b1001111010001,
13'b1001111100000,
13'b1010110000000,
13'b1010110000001,
13'b1010110010000,
13'b1010110010001,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010111000000,
13'b1010111000001,
13'b1010111010000,
13'b1011110010000,
13'b1011110100000,
13'b1011110100001,
13'b1011110110000,
13'b1011110110001,
13'b1011111000000: edge_mask_reg_512p3[411] <= 1'b1;
 		default: edge_mask_reg_512p3[411] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010110,
13'b1010010111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000110,
13'b101010000111,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000110,
13'b110010000111,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000110110,
13'b111000110111,
13'b111001000110,
13'b111001000111,
13'b111001010110,
13'b111001010111,
13'b1000000010110,
13'b1000000010111,
13'b1000000011000,
13'b1000000100110,
13'b1000000100111,
13'b1000000110110,
13'b1000000110111,
13'b1000001000110,
13'b1000001000111,
13'b1000001010110,
13'b1000001010111,
13'b1001000010110,
13'b1001000010111,
13'b1001000011000,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110110,
13'b1001000110111,
13'b1001001000110,
13'b1001001000111,
13'b1001001010110,
13'b1001001010111,
13'b1010000000110,
13'b1010000000111,
13'b1010000001000,
13'b1010000010110,
13'b1010000010111,
13'b1010000011000,
13'b1010000100110,
13'b1010000100111,
13'b1010000101000,
13'b1010000110110,
13'b1010000110111,
13'b1010001000110,
13'b1010001000111,
13'b1010001010110,
13'b1010001010111,
13'b1011000000110,
13'b1011000000111,
13'b1011000001000,
13'b1011000010110,
13'b1011000010111,
13'b1011000011000,
13'b1011000100110,
13'b1011000100111,
13'b1011000101000,
13'b1011000110110,
13'b1011000110111,
13'b1011001000110,
13'b1011001000111,
13'b1011001010110,
13'b1011001010111,
13'b1100000000110,
13'b1100000000111,
13'b1100000010110,
13'b1100000010111,
13'b1100000011000,
13'b1100000100110,
13'b1100000100111,
13'b1100000101000,
13'b1100000110110,
13'b1100000110111,
13'b1100001000110,
13'b1100001000111,
13'b1100001010110,
13'b1100001010111,
13'b1101000000100,
13'b1101000000101,
13'b1101000000110,
13'b1101000000111,
13'b1101000001000,
13'b1101000010100,
13'b1101000010101,
13'b1101000010110,
13'b1101000010111,
13'b1101000011000,
13'b1101000100100,
13'b1101000100101,
13'b1101000100110,
13'b1101000100111,
13'b1101000101000,
13'b1101000110100,
13'b1101000110101,
13'b1101000110110,
13'b1101000110111,
13'b1101000111000,
13'b1101001000100,
13'b1101001000101,
13'b1101001000110,
13'b1101001000111,
13'b1101001001000,
13'b1101001010110,
13'b1101001010111,
13'b1110000000100,
13'b1110000000101,
13'b1110000000110,
13'b1110000000111,
13'b1110000001000,
13'b1110000010100,
13'b1110000010101,
13'b1110000010110,
13'b1110000010111,
13'b1110000011000,
13'b1110000100100,
13'b1110000100101,
13'b1110000100110,
13'b1110000100111,
13'b1110000101000,
13'b1110000110100,
13'b1110000110101,
13'b1110000110110,
13'b1110000110111,
13'b1110000111000,
13'b1110001000100,
13'b1110001000101,
13'b1110001000110,
13'b1110001000111,
13'b1110001001000,
13'b1110001010100,
13'b1110001010101,
13'b1110001010110,
13'b1110001010111,
13'b1111000000100,
13'b1111000000101,
13'b1111000000110,
13'b1111000000111,
13'b1111000001000,
13'b1111000010100,
13'b1111000010101,
13'b1111000010110,
13'b1111000010111,
13'b1111000011000,
13'b1111000100100,
13'b1111000100101,
13'b1111000100110,
13'b1111000100111,
13'b1111000101000,
13'b1111000110100,
13'b1111000110101,
13'b1111000110110,
13'b1111000110111,
13'b1111000111000,
13'b1111001000100,
13'b1111001000101,
13'b1111001000110,
13'b1111001000111,
13'b1111001010110,
13'b1111001010111: edge_mask_reg_512p3[412] <= 1'b1;
 		default: edge_mask_reg_512p3[412] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b10001111010,
13'b10001111011,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b11001111010,
13'b11001111011,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011011100,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011101100,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b111010111000,
13'b111010111001,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b1000010111000,
13'b1000010111001,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011101001,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001011111001,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1011010110111,
13'b1011010111000,
13'b1011010111001,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011001001,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011011001,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011101000,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011011111000,
13'b1011100000110,
13'b1011100000111,
13'b1011100001000,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100011111000,
13'b1100100000110,
13'b1100100000111,
13'b1100100001000,
13'b1101011000101,
13'b1101011000110,
13'b1101011000111,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011100100,
13'b1101011100101,
13'b1101011100110,
13'b1101011100111,
13'b1101011110100,
13'b1101011110101,
13'b1101011110110,
13'b1101011110111,
13'b1110011000110,
13'b1110011010101,
13'b1110011010110,
13'b1110011100101,
13'b1110011100110,
13'b1110011110101,
13'b1110011110110,
13'b1111011010101,
13'b1111011010110,
13'b1111011100101,
13'b1111011100110,
13'b1111011110101: edge_mask_reg_512p3[413] <= 1'b1;
 		default: edge_mask_reg_512p3[413] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101011000,
13'b101011001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001001,
13'b10101001010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001001,
13'b11101001010,
13'b100001111000,
13'b100001111001,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111001,
13'b100100111010,
13'b100101001001,
13'b100101001010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b110010001000,
13'b110010001001,
13'b110010011000,
13'b110010011001,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b111010100110,
13'b111010100111,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b1000010100110,
13'b1000010100111,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011101001,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001011111001,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1010010100101,
13'b1010010100110,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110010,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011101000,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011011111000,
13'b1011100000110,
13'b1011100000111,
13'b1011100001000,
13'b1100010100010,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100011000010,
13'b1100011000011,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010011,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100011,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100011111000,
13'b1100100000110,
13'b1100100000111,
13'b1100100001000,
13'b1101010110011,
13'b1101010110100,
13'b1101010110101,
13'b1101010110110,
13'b1101011000010,
13'b1101011000011,
13'b1101011000100,
13'b1101011000101,
13'b1101011000110,
13'b1101011000111,
13'b1101011010011,
13'b1101011010100,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011100011,
13'b1101011100100,
13'b1101011100101,
13'b1101011100110,
13'b1101011100111,
13'b1101011110100,
13'b1101011110101,
13'b1101011110110,
13'b1101011110111,
13'b1110010110011,
13'b1110011000011,
13'b1110011000100,
13'b1110011000101,
13'b1110011010011,
13'b1110011010100,
13'b1110011010101,
13'b1110011010110,
13'b1110011100011,
13'b1110011100100,
13'b1110011100101,
13'b1110011100110,
13'b1110011110100,
13'b1110011110101,
13'b1110011110110,
13'b1111011010100,
13'b1111011010101,
13'b1111011100101,
13'b1111011100110,
13'b1111011110101: edge_mask_reg_512p3[414] <= 1'b1;
 		default: edge_mask_reg_512p3[414] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110001,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000000,
13'b11110000001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010000,
13'b11110010001,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100000,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110000,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100100111,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010000,
13'b100110010001,
13'b100110010010,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100000,
13'b100110100001,
13'b100110100100,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110000,
13'b100110110001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000000,
13'b100111000001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100100111,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100000,
13'b101110100001,
13'b101110100010,
13'b101110100011,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110000,
13'b101110110001,
13'b101110110010,
13'b101110110011,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000000,
13'b101111000001,
13'b101111000010,
13'b101111000100,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010000,
13'b101111010001,
13'b101111010010,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110011,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000000,
13'b110111000001,
13'b110111000010,
13'b110111000011,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010000,
13'b110111010001,
13'b110111010010,
13'b110111010011,
13'b110111010100,
13'b110111010101,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100111,
13'b111101101000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110111,
13'b111101111000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110111000,
13'b111111000000,
13'b111111000001,
13'b111111000010,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111010000,
13'b111111010001,
13'b111111010010,
13'b111111010011,
13'b111111010100,
13'b111111010101,
13'b1000101100001,
13'b1000101100010,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111010010,
13'b1000111010011,
13'b1000111010100,
13'b1001110000010,
13'b1001110010010,
13'b1001110010011,
13'b1001110100010,
13'b1001110100011,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100: edge_mask_reg_512p3[415] <= 1'b1;
 		default: edge_mask_reg_512p3[415] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110001,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000000,
13'b11110000001,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010000,
13'b11110010001,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100000,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110000,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100100111,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110000,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000000,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010000,
13'b100110010001,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100000,
13'b100110100001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110000,
13'b100110110001,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b101100100111,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110000,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000000,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010000,
13'b101110010001,
13'b101110010010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100000,
13'b101110100001,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110000,
13'b101110110001,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111001001,
13'b101111010111,
13'b101111011000,
13'b101111011001,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110000,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000000,
13'b110110000001,
13'b110110000010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010000,
13'b110110010001,
13'b110110010010,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110100000,
13'b110110100001,
13'b110110100010,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110110000,
13'b110110110001,
13'b110110110010,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110110111010,
13'b110111000111,
13'b110111001000,
13'b110111001001,
13'b110111010111,
13'b110111011000,
13'b110111011001,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101100001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100111,
13'b111101101000,
13'b111101110001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000000,
13'b111110000001,
13'b111110000010,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110010000,
13'b111110010001,
13'b111110010010,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110100000,
13'b111110100001,
13'b111110100010,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110101001,
13'b111110110000,
13'b111110110001,
13'b111110110010,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111111000001,
13'b111111000010,
13'b111111000101,
13'b111111000110,
13'b1000101010010,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110010111,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110100111,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000110110111,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000101,
13'b1000111000110,
13'b1001101100010,
13'b1001101100011,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110100110,
13'b1001110100111,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001110110110,
13'b1001110110111,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111000110,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110010101,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110100101,
13'b1010110100110,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010110110101,
13'b1010110110110,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111000101,
13'b1011110000011,
13'b1011110000100,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110010101,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110100101,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011110110100,
13'b1011110110101,
13'b1011111000010,
13'b1011111000011,
13'b1011111000100,
13'b1100110010100,
13'b1100110100011,
13'b1100110100100,
13'b1100110100101,
13'b1100110110011,
13'b1100110110100,
13'b1100110110101: edge_mask_reg_512p3[416] <= 1'b1;
 		default: edge_mask_reg_512p3[416] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000110111,
13'b100000111000,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110111,
13'b101000111000,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b1000000010010,
13'b1000000010011,
13'b1010000000010,
13'b1010000000011: edge_mask_reg_512p3[417] <= 1'b1;
 		default: edge_mask_reg_512p3[417] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000110111,
13'b100000111000,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b110000100111,
13'b110000101000,
13'b1010000000010,
13'b1010000000011: edge_mask_reg_512p3[418] <= 1'b1;
 		default: edge_mask_reg_512p3[418] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[419] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[420] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[421] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b10001101001,
13'b10001101010,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010011,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100011,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110010,
13'b10010110011,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000010,
13'b10011000011,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000101,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010011,
13'b101010010100,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111001,
13'b101100111010,
13'b101101001001,
13'b101101001010,
13'b110010100001,
13'b110010100010,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010111001,
13'b110010111010,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011001001,
13'b110011001010,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011001,
13'b110011011010,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101001,
13'b110011101010,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111001,
13'b110011111010,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b111010110001,
13'b111010110010,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b1000011010010,
13'b1000011010011,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110100,
13'b1000100110101,
13'b1001011100010,
13'b1001011100011,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1010011110010,
13'b1010011110011,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010010,
13'b1010100010011,
13'b1010100100010,
13'b1010100100011: edge_mask_reg_512p3[422] <= 1'b1;
 		default: edge_mask_reg_512p3[422] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111010,
13'b10001101001,
13'b10001101010,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010011,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100011,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110010,
13'b10010110011,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000010,
13'b10011000011,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b10101111011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000101,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011010001,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011100010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110001,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000010,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111001,
13'b101100111010,
13'b101101000100,
13'b101101000101,
13'b110010110001,
13'b110010110010,
13'b110010111001,
13'b110010111010,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011001001,
13'b110011001010,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011011001,
13'b110011011010,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011101001,
13'b110011101010,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011111001,
13'b110011111010,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100110100,
13'b110100110101,
13'b111011100010,
13'b111011100011,
13'b111011110010,
13'b111011110011,
13'b111100000010,
13'b111100000011,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100100010,
13'b111100100011,
13'b1000100010011: edge_mask_reg_512p3[423] <= 1'b1;
 		default: edge_mask_reg_512p3[423] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b11110111100,
13'b100100111001,
13'b100100111010,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b100111001000,
13'b100111001001,
13'b100111001010,
13'b100111001011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110011011,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110101011,
13'b101110111000,
13'b101110111001,
13'b101110111010,
13'b101110111011,
13'b101111001000,
13'b101111001001,
13'b101111001010,
13'b101111001011,
13'b101111011001,
13'b101111011010,
13'b110101101000,
13'b110101101001,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110001011,
13'b110110011000,
13'b110110011001,
13'b110110011010,
13'b110110011011,
13'b110110101000,
13'b110110101001,
13'b110110101010,
13'b110110101011,
13'b110110111001,
13'b110110111010,
13'b110110111011,
13'b110111001010,
13'b110111001011,
13'b111101111000,
13'b111101111001,
13'b111101111010,
13'b111110000111,
13'b111110001000,
13'b111110001001,
13'b111110001010,
13'b111110001011,
13'b111110010111,
13'b111110011000,
13'b111110011001,
13'b111110011010,
13'b111110011011,
13'b111110101000,
13'b111110101001,
13'b111110101010,
13'b111110101011,
13'b111110111001,
13'b111110111010,
13'b111110111011,
13'b111111001010,
13'b111111001011,
13'b1000101101000,
13'b1000101111000,
13'b1000101111001,
13'b1000101111010,
13'b1000110000111,
13'b1000110001000,
13'b1000110001001,
13'b1000110001010,
13'b1000110001011,
13'b1000110010111,
13'b1000110011000,
13'b1000110011001,
13'b1000110011010,
13'b1000110011011,
13'b1000110101000,
13'b1000110101001,
13'b1000110101010,
13'b1000110101011,
13'b1000110111001,
13'b1000110111010,
13'b1000110111011,
13'b1000111001010,
13'b1000111001011,
13'b1001101101000,
13'b1001101110111,
13'b1001101111000,
13'b1001101111001,
13'b1001101111010,
13'b1001110000111,
13'b1001110001000,
13'b1001110001001,
13'b1001110001010,
13'b1001110001011,
13'b1001110010111,
13'b1001110011000,
13'b1001110011001,
13'b1001110011010,
13'b1001110011011,
13'b1001110011100,
13'b1001110101000,
13'b1001110101001,
13'b1001110101010,
13'b1001110101011,
13'b1001110111001,
13'b1001110111010,
13'b1001110111011,
13'b1001111001010,
13'b1001111001011,
13'b1010101101000,
13'b1010101111000,
13'b1010101111001,
13'b1010101111010,
13'b1010110000111,
13'b1010110001000,
13'b1010110001001,
13'b1010110001010,
13'b1010110001011,
13'b1010110010111,
13'b1010110011000,
13'b1010110011001,
13'b1010110011010,
13'b1010110011011,
13'b1010110100111,
13'b1010110101000,
13'b1010110101001,
13'b1010110101010,
13'b1010110101011,
13'b1010110111001,
13'b1010110111010,
13'b1010110111011,
13'b1010111001010,
13'b1010111001011,
13'b1011101101000,
13'b1011101101001,
13'b1011101110111,
13'b1011101111000,
13'b1011101111001,
13'b1011101111010,
13'b1011110000111,
13'b1011110001000,
13'b1011110001001,
13'b1011110001010,
13'b1011110001011,
13'b1011110010111,
13'b1011110011000,
13'b1011110011001,
13'b1011110011010,
13'b1011110011011,
13'b1011110011100,
13'b1011110100111,
13'b1011110101000,
13'b1011110101001,
13'b1011110101010,
13'b1011110101011,
13'b1011110101100,
13'b1011110111000,
13'b1011110111001,
13'b1011110111010,
13'b1011110111011,
13'b1011111001010,
13'b1011111001011,
13'b1100101101000,
13'b1100101110111,
13'b1100101111000,
13'b1100101111001,
13'b1100101111010,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1100110001001,
13'b1100110001010,
13'b1100110001011,
13'b1100110010110,
13'b1100110010111,
13'b1100110011000,
13'b1100110011001,
13'b1100110011010,
13'b1100110011011,
13'b1100110011100,
13'b1100110100111,
13'b1100110101000,
13'b1100110101001,
13'b1100110101010,
13'b1100110101011,
13'b1100110101100,
13'b1100110111000,
13'b1100110111001,
13'b1100110111010,
13'b1100110111011,
13'b1100111001010,
13'b1100111001011,
13'b1101101101000,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101101111001,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1101110001001,
13'b1101110001010,
13'b1101110001011,
13'b1101110010110,
13'b1101110010111,
13'b1101110011000,
13'b1101110011001,
13'b1101110011010,
13'b1101110011011,
13'b1101110100111,
13'b1101110101000,
13'b1101110101001,
13'b1101110101010,
13'b1101110101011,
13'b1101110111000,
13'b1101110111001,
13'b1101110111010,
13'b1101110111011,
13'b1101111001010,
13'b1101111001011,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110101111001,
13'b1110110000110,
13'b1110110000111,
13'b1110110001000,
13'b1110110001001,
13'b1110110001010,
13'b1110110010110,
13'b1110110010111,
13'b1110110011000,
13'b1110110011001,
13'b1110110011010,
13'b1110110011011,
13'b1110110100111,
13'b1110110101000,
13'b1110110101001,
13'b1110110101010,
13'b1110110101011,
13'b1110110111010,
13'b1111101110110,
13'b1111101110111,
13'b1111101111000,
13'b1111110000110,
13'b1111110000111,
13'b1111110001000,
13'b1111110001001,
13'b1111110001010,
13'b1111110010110,
13'b1111110010111,
13'b1111110011000,
13'b1111110011001,
13'b1111110011010,
13'b1111110011011,
13'b1111110101000,
13'b1111110101001,
13'b1111110101010,
13'b1111110101011,
13'b1111110111010: edge_mask_reg_512p3[424] <= 1'b1;
 		default: edge_mask_reg_512p3[424] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010101,
13'b11101010110,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101010101,
13'b100101010110,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101010101,
13'b101101010110,
13'b110001100110,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110101000101,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100010,
13'b1000100100011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100010,
13'b1001100100011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100100010,
13'b1010100100011,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011100101,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011011110101,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1100010010100,
13'b1100010010101,
13'b1100010010110,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100011000010,
13'b1100011000011,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011010001,
13'b1100011010010,
13'b1100011010011,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011100000,
13'b1100011100001,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011100101,
13'b1100011110000,
13'b1100011110001,
13'b1100011110010,
13'b1100011110011,
13'b1100011110100,
13'b1100100000000,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100000100,
13'b1100100010000,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100100001,
13'b1100100100010,
13'b1101010010100,
13'b1101010010101,
13'b1101010010110,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010100110,
13'b1101010110010,
13'b1101010110011,
13'b1101010110100,
13'b1101010110101,
13'b1101010110110,
13'b1101011000010,
13'b1101011000011,
13'b1101011000100,
13'b1101011000101,
13'b1101011000110,
13'b1101011010001,
13'b1101011010010,
13'b1101011010011,
13'b1101011010100,
13'b1101011010101,
13'b1101011100000,
13'b1101011100001,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011100101,
13'b1101011110000,
13'b1101011110001,
13'b1101011110010,
13'b1101011110011,
13'b1101011110100,
13'b1101100000000,
13'b1101100000001,
13'b1101100000010,
13'b1101100000011,
13'b1101100000100,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100100001,
13'b1101100100010,
13'b1110010010100,
13'b1110010010101,
13'b1110010010110,
13'b1110010100011,
13'b1110010100100,
13'b1110010100101,
13'b1110010100110,
13'b1110010110010,
13'b1110010110011,
13'b1110010110100,
13'b1110010110101,
13'b1110010110110,
13'b1110011000001,
13'b1110011000010,
13'b1110011000011,
13'b1110011000100,
13'b1110011000101,
13'b1110011000110,
13'b1110011010000,
13'b1110011010001,
13'b1110011010010,
13'b1110011010011,
13'b1110011010100,
13'b1110011010101,
13'b1110011100000,
13'b1110011100001,
13'b1110011100010,
13'b1110011100011,
13'b1110011100100,
13'b1110011100101,
13'b1110011110000,
13'b1110011110001,
13'b1110011110010,
13'b1110011110011,
13'b1110011110100,
13'b1110100000000,
13'b1110100000001,
13'b1110100000010,
13'b1110100000011,
13'b1110100010000,
13'b1110100010001,
13'b1111010010100,
13'b1111010010101,
13'b1111010100011,
13'b1111010100100,
13'b1111010100101,
13'b1111010100110,
13'b1111010110010,
13'b1111010110011,
13'b1111010110100,
13'b1111010110101,
13'b1111010110110,
13'b1111011000001,
13'b1111011000010,
13'b1111011000011,
13'b1111011000100,
13'b1111011000101,
13'b1111011000110,
13'b1111011010000,
13'b1111011010001,
13'b1111011010010,
13'b1111011010011,
13'b1111011010100,
13'b1111011010101,
13'b1111011100000,
13'b1111011100001,
13'b1111011100010,
13'b1111011100011,
13'b1111011100100,
13'b1111011110000,
13'b1111011110001,
13'b1111011110010,
13'b1111100000000,
13'b1111100000001: edge_mask_reg_512p3[425] <= 1'b1;
 		default: edge_mask_reg_512p3[425] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011110110,
13'b11011110111,
13'b100001000101,
13'b100001000110,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011110110,
13'b100011110111,
13'b101001000101,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011110110,
13'b101011110111,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b111001110100,
13'b111001110101,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000101,
13'b1000011000110,
13'b1001001110100,
13'b1001001110101,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1010001110100,
13'b1010001110101,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000101,
13'b1011001110100,
13'b1011001110101,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000101,
13'b1011011000110,
13'b1100001110011,
13'b1100001110100,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010010110,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100011000101,
13'b1100011000110,
13'b1101001110011,
13'b1101001110100,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010010101,
13'b1101010010110,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010100110,
13'b1101010110011,
13'b1101010110100,
13'b1101010110101,
13'b1101010110110,
13'b1101011000101,
13'b1101011000110,
13'b1110001110011,
13'b1110001110100,
13'b1110010000010,
13'b1110010000011,
13'b1110010000100,
13'b1110010000101,
13'b1110010010001,
13'b1110010010010,
13'b1110010010011,
13'b1110010010100,
13'b1110010010101,
13'b1110010010110,
13'b1110010100010,
13'b1110010100011,
13'b1110010100100,
13'b1110010100101,
13'b1110010100110,
13'b1110010110011,
13'b1110010110100,
13'b1110010110101,
13'b1110010110110,
13'b1110011000101,
13'b1110011000110,
13'b1111010000010,
13'b1111010000011,
13'b1111010000100,
13'b1111010000101,
13'b1111010010001,
13'b1111010010010,
13'b1111010010011,
13'b1111010010100,
13'b1111010010101,
13'b1111010100001,
13'b1111010100010,
13'b1111010100011,
13'b1111010100100,
13'b1111010100101,
13'b1111010100110,
13'b1111010110010,
13'b1111010110011,
13'b1111010110100,
13'b1111010110101,
13'b1111010110110,
13'b1111011000100,
13'b1111011000101: edge_mask_reg_512p3[426] <= 1'b1;
 		default: edge_mask_reg_512p3[426] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000100,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b11001000011,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010101,
13'b11010010110,
13'b100000110010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000001,
13'b100001000010,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010001,
13'b100001010010,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100001,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010010101,
13'b100010010110,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000000,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010000,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100000,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000101,
13'b101010000110,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110000,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010000,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100000,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110010000101,
13'b110010000110,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010101,
13'b111001010110,
13'b111001100000,
13'b111001100001,
13'b111001100010,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001100000,
13'b1000001100001,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001010000,
13'b1001001010001,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000110000,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1101000100000,
13'b1101000100001,
13'b1110000000000,
13'b1110000000001,
13'b1110000000010,
13'b1110000010000,
13'b1110000010001,
13'b1110000100000,
13'b1111000000000,
13'b1111000000001,
13'b1111000010000,
13'b1111000010001: edge_mask_reg_512p3[427] <= 1'b1;
 		default: edge_mask_reg_512p3[427] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010110,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000110,
13'b110001000111,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100001,
13'b1000000100010,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000100010,
13'b1100000100011,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1110000000000,
13'b1110000000001,
13'b1110000000010,
13'b1110000010000,
13'b1110000010001,
13'b1111000000000,
13'b1111000000001,
13'b1111000010000,
13'b1111000010001: edge_mask_reg_512p3[428] <= 1'b1;
 		default: edge_mask_reg_512p3[428] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010101,
13'b11010010110,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010101,
13'b100010010110,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000101,
13'b101010000110,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000101,
13'b110010000110,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001100000,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001010000,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001100000,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001100000,
13'b1010001100001,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001010000,
13'b1011001010001,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100001000000,
13'b1100001010000,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1101000100000,
13'b1101000100001,
13'b1101000110000,
13'b1101000110001,
13'b1101001000000,
13'b1110000000000,
13'b1110000000001,
13'b1110000000010,
13'b1110000010000,
13'b1110000010001,
13'b1110000100000,
13'b1110000100001,
13'b1110000110000,
13'b1111000000000,
13'b1111000000001,
13'b1111000010000,
13'b1111000010001: edge_mask_reg_512p3[429] <= 1'b1;
 		default: edge_mask_reg_512p3[429] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101010,
13'b10110101011,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110011010,
13'b11110011011,
13'b11110101011,
13'b100010111001,
13'b100010111010,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111010,
13'b100101111011,
13'b101011001001,
13'b101011001010,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101101000,
13'b101101101001,
13'b110011010110,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101100111,
13'b1000101101000,
13'b1001011100101,
13'b1001011100110,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100101000,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101100110,
13'b1001101100111,
13'b1010011100101,
13'b1010011100110,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1011011110011,
13'b1011011110100,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1100100000011,
13'b1100100000100,
13'b1100100010011,
13'b1100100010100,
13'b1100100010101,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100110100,
13'b1100100110101,
13'b1100100110110,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1101100100101,
13'b1101100110101,
13'b1101100110110,
13'b1101101000101,
13'b1101101000110,
13'b1101101010110: edge_mask_reg_512p3[430] <= 1'b1;
 		default: edge_mask_reg_512p3[430] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001010,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b1011011011,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10011101010,
13'b10011101011,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111010,
13'b11110111011,
13'b100100001011,
13'b100100011011,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110001001,
13'b110100101000,
13'b110100101001,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110001000,
13'b110110001001,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110001000,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101101001,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000111,
13'b1001100100111,
13'b1001100101000,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000111,
13'b1010100100111,
13'b1010100101000,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101010101,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101110111,
13'b1010101111000,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000101,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010101,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100101,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1100100110101,
13'b1100100110110,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101100101,
13'b1100101100110,
13'b1100101100111,
13'b1101100110110,
13'b1101101000110,
13'b1101101010110,
13'b1101101100110: edge_mask_reg_512p3[431] <= 1'b1;
 		default: edge_mask_reg_512p3[431] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[432] <= 1'b0;
 	endcase

    case({x,y,z})
13'b101000100100,
13'b101000100101: edge_mask_reg_512p3[433] <= 1'b1;
 		default: edge_mask_reg_512p3[433] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010101000,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000111,
13'b110110001000,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b1000011100110,
13'b1000011100111,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100001000,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100011000,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1001011100101,
13'b1001011100110,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100010111,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1010011100101,
13'b1010011100110,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100000111,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1010100010111,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1011011100101,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1100011100101,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1100100000011,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100010101,
13'b1100100010110,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100100110101,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101000101,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1101011110011,
13'b1101011110100,
13'b1101011110101,
13'b1101100000010,
13'b1101100000011,
13'b1101100000100,
13'b1101100000101,
13'b1101100000110,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100010100,
13'b1101100010101,
13'b1101100010110,
13'b1101100100001,
13'b1101100100010,
13'b1101100100011,
13'b1101100100100,
13'b1101100100101,
13'b1101100100110,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101100110100,
13'b1101100110101,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101000100,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1110100000010,
13'b1110100000011,
13'b1110100000100,
13'b1110100010010,
13'b1110100010011,
13'b1110100010100,
13'b1110100100001,
13'b1110100100010,
13'b1110100100011,
13'b1110100110001,
13'b1110100110010,
13'b1110100110011,
13'b1110101000001,
13'b1110101000010,
13'b1110101010001,
13'b1111100000011,
13'b1111100000100,
13'b1111100010010,
13'b1111100010011,
13'b1111100010100,
13'b1111100100010,
13'b1111100100011: edge_mask_reg_512p3[434] <= 1'b1;
 		default: edge_mask_reg_512p3[434] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010010110,
13'b1010010111,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b101010100110,
13'b101010100111,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000111,
13'b110110001000,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b1000011000010,
13'b1000011000011,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1001011000001,
13'b1001011000010,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1011011010000,
13'b1011011010001,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011100000000,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100100000,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1100011010000,
13'b1100011100000,
13'b1100011100001,
13'b1100011110000,
13'b1100011110001,
13'b1100100000000,
13'b1100100000001,
13'b1100100000010,
13'b1100100010000,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100100000,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1101011100000,
13'b1101011110000,
13'b1101011110001,
13'b1101100000000,
13'b1101100000001,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100100000,
13'b1101100100001,
13'b1101100100010,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101000100,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1110100010001,
13'b1110100100001,
13'b1110100110001,
13'b1110100110010,
13'b1110101000001,
13'b1110101010001: edge_mask_reg_512p3[435] <= 1'b1;
 		default: edge_mask_reg_512p3[435] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110010,
13'b110011110011,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000111,
13'b110110001000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000111,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1001011110001,
13'b1001011110010,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1010100000010,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1011100010000,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100100000,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1100100100000,
13'b1100100100001,
13'b1100100100010,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1101100100000,
13'b1101100100001,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101000100,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1110100110001,
13'b1110100110010,
13'b1110101000001,
13'b1110101010001: edge_mask_reg_512p3[436] <= 1'b1;
 		default: edge_mask_reg_512p3[436] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10011000110,
13'b10011000111,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b101011010110,
13'b101011010111,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000111,
13'b110110001000,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b1000011110100,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1001011110100,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100010001,
13'b1011100010010,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100100001,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1100100000001,
13'b1100100000010,
13'b1100100000011,
13'b1100100010001,
13'b1100100010010,
13'b1100100010011,
13'b1100100010100,
13'b1100100100000,
13'b1100100100001,
13'b1100100100010,
13'b1100100100011,
13'b1100100100100,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1101100000001,
13'b1101100000010,
13'b1101100010000,
13'b1101100010001,
13'b1101100010010,
13'b1101100010011,
13'b1101100100000,
13'b1101100100001,
13'b1101100100010,
13'b1101100100011,
13'b1101100100100,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101100110100,
13'b1101101000000,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101000100,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1110100000000,
13'b1110100000001,
13'b1110100010000,
13'b1110100010001,
13'b1110100010010,
13'b1110100100000,
13'b1110100100001,
13'b1110100100010,
13'b1110100110000,
13'b1110100110001,
13'b1110100110010,
13'b1110101000001,
13'b1110101000010,
13'b1110101010001,
13'b1111100010001,
13'b1111100010010,
13'b1111100100001,
13'b1111100100010,
13'b1111100110001: edge_mask_reg_512p3[437] <= 1'b1;
 		default: edge_mask_reg_512p3[437] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b100011101000,
13'b100011101001,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b101011101000,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b110011111000,
13'b110011111001,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000111,
13'b110110001000,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100010111,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100100111,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100100110,
13'b1001100100111,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001100110111,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101000111,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100100101,
13'b1010100100110,
13'b1010100100111,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010100110110,
13'b1010100110111,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101000110,
13'b1010101000111,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1011100100010,
13'b1011100100011,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101000110,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1100100100011,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100110000,
13'b1100100110001,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100100110101,
13'b1100100110110,
13'b1100101000000,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101000101,
13'b1100101000110,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101010101,
13'b1101100100011,
13'b1101100100100,
13'b1101100100101,
13'b1101100110000,
13'b1101100110001,
13'b1101100110010,
13'b1101100110011,
13'b1101100110100,
13'b1101100110101,
13'b1101100110110,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101000100,
13'b1101101000101,
13'b1101101000110,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101010100,
13'b1110100100011,
13'b1110100100100,
13'b1110100110001,
13'b1110100110010,
13'b1110100110011,
13'b1110100110100,
13'b1110101000001,
13'b1110101000010,
13'b1110101000011,
13'b1110101000100,
13'b1110101010001,
13'b1110101010010,
13'b1111100110011,
13'b1111101000010,
13'b1111101000011,
13'b1111101000100: edge_mask_reg_512p3[438] <= 1'b1;
 		default: edge_mask_reg_512p3[438] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[439] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101011,
13'b10101100,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b10111101,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11001101,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11011101,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11101101,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b11111101,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100001101,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100011101,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100101101,
13'b100111010,
13'b100111011,
13'b100111100,
13'b100111101,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101001101,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101011101,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b101101101,
13'b1010111011,
13'b1010111100,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011011101,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011101101,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1011111101,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100001101,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100011101,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100101101,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1100111101,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101001101,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101011101,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101101101,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1101111101,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110001101,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b1110011101,
13'b10011001011,
13'b10011001100,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100011101,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100101101,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10100111101,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101001101,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101011101,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101101101,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001011,
13'b10110001100,
13'b10110011011,
13'b10110011100,
13'b11011101011,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100011101,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100101101,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11100111101,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101001101,
13'b11101001110,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101011101,
13'b11101011110,
13'b11101101100,
13'b11101101101,
13'b100100001010,
13'b100100001011,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100011101,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100101101,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100100111101,
13'b100100111110,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101001101,
13'b100101001110,
13'b100101011011,
13'b100101011100,
13'b100101011101,
13'b100101011110,
13'b100101101100,
13'b100101101101,
13'b101100001010,
13'b101100001011,
13'b101100001100,
13'b101100011010,
13'b101100011011,
13'b101100011100,
13'b101100011101,
13'b101100101010,
13'b101100101011,
13'b101100101100,
13'b101100101101,
13'b101100111010,
13'b101100111011,
13'b101100111100,
13'b101100111101,
13'b101100111110,
13'b101101001010,
13'b101101001011,
13'b101101001100,
13'b101101001101,
13'b101101001110,
13'b101101011010,
13'b101101011011,
13'b101101011100,
13'b101101011101,
13'b101101011110,
13'b101101101100,
13'b101101101101,
13'b110100001010,
13'b110100001011,
13'b110100001100,
13'b110100011001,
13'b110100011010,
13'b110100011011,
13'b110100011100,
13'b110100011101,
13'b110100011110,
13'b110100101001,
13'b110100101010,
13'b110100101011,
13'b110100101100,
13'b110100101101,
13'b110100101110,
13'b110100111010,
13'b110100111011,
13'b110100111100,
13'b110100111101,
13'b110100111110,
13'b110101001010,
13'b110101001011,
13'b110101001100,
13'b110101001101,
13'b110101001110,
13'b110101011010,
13'b110101011011,
13'b110101011100,
13'b110101011101,
13'b110101011110,
13'b110101101100,
13'b110101101101,
13'b111100001010,
13'b111100001011,
13'b111100001100,
13'b111100011001,
13'b111100011010,
13'b111100011011,
13'b111100011100,
13'b111100011101,
13'b111100011110,
13'b111100101001,
13'b111100101010,
13'b111100101011,
13'b111100101100,
13'b111100101101,
13'b111100101110,
13'b111100111010,
13'b111100111011,
13'b111100111100,
13'b111100111101,
13'b111100111110,
13'b111101001001,
13'b111101001010,
13'b111101001011,
13'b111101001100,
13'b111101001101,
13'b111101001110,
13'b111101011010,
13'b111101011011,
13'b111101011100,
13'b111101011101,
13'b111101011110,
13'b111101101101,
13'b111101101110,
13'b1000100001010,
13'b1000100001011,
13'b1000100011001,
13'b1000100011010,
13'b1000100011011,
13'b1000100011100,
13'b1000100011101,
13'b1000100011110,
13'b1000100101001,
13'b1000100101010,
13'b1000100101011,
13'b1000100101100,
13'b1000100101101,
13'b1000100101110,
13'b1000100111001,
13'b1000100111010,
13'b1000100111011,
13'b1000100111100,
13'b1000100111101,
13'b1000100111110,
13'b1000101001001,
13'b1000101001010,
13'b1000101001011,
13'b1000101001100,
13'b1000101001101,
13'b1000101001110,
13'b1000101011011,
13'b1000101011100,
13'b1000101011101,
13'b1000101011110,
13'b1000101101101,
13'b1001100001001,
13'b1001100001010,
13'b1001100001011,
13'b1001100011001,
13'b1001100011010,
13'b1001100011011,
13'b1001100011100,
13'b1001100011101,
13'b1001100011110,
13'b1001100101001,
13'b1001100101010,
13'b1001100101011,
13'b1001100101100,
13'b1001100101101,
13'b1001100101110,
13'b1001100111001,
13'b1001100111010,
13'b1001100111011,
13'b1001100111100,
13'b1001100111101,
13'b1001100111110,
13'b1001101001001,
13'b1001101001010,
13'b1001101001011,
13'b1001101001100,
13'b1001101001101,
13'b1001101001110,
13'b1001101011010,
13'b1001101011011,
13'b1001101011100,
13'b1001101011101,
13'b1001101011110,
13'b1001101101101,
13'b1010100001001,
13'b1010100001010,
13'b1010100001011,
13'b1010100011001,
13'b1010100011010,
13'b1010100011011,
13'b1010100011100,
13'b1010100011101,
13'b1010100101000,
13'b1010100101001,
13'b1010100101010,
13'b1010100101011,
13'b1010100101100,
13'b1010100101101,
13'b1010100111000,
13'b1010100111001,
13'b1010100111010,
13'b1010100111011,
13'b1010100111100,
13'b1010100111101,
13'b1010100111110,
13'b1010101001001,
13'b1010101001010,
13'b1010101001011,
13'b1010101001100,
13'b1010101001101,
13'b1010101001110,
13'b1010101011010,
13'b1010101011011,
13'b1010101011100,
13'b1010101011101,
13'b1011100001010,
13'b1011100011001,
13'b1011100011010,
13'b1011100011011,
13'b1011100101000,
13'b1011100101001,
13'b1011100101010,
13'b1011100101011,
13'b1011100101100,
13'b1011100101101,
13'b1011100111000,
13'b1011100111001,
13'b1011100111010,
13'b1011100111011,
13'b1011100111100,
13'b1011100111101,
13'b1011100111110,
13'b1011101001001,
13'b1011101001010,
13'b1011101001011,
13'b1011101001100,
13'b1011101001101,
13'b1011101001110,
13'b1011101011100,
13'b1011101011101,
13'b1100100011000,
13'b1100100011001,
13'b1100100100111,
13'b1100100101000,
13'b1100100101001,
13'b1100100101010,
13'b1100100101011,
13'b1100100101100,
13'b1100100110111,
13'b1100100111000,
13'b1100100111001,
13'b1100100111010,
13'b1100100111011,
13'b1100100111100,
13'b1100100111101,
13'b1100100111110,
13'b1100101001000,
13'b1100101001001,
13'b1100101001010,
13'b1100101001011,
13'b1100101001100,
13'b1100101001101,
13'b1100101001110,
13'b1100101011100,
13'b1100101011101,
13'b1101100011000,
13'b1101100101000,
13'b1101100101001,
13'b1101100101010,
13'b1101100101011,
13'b1101100111000,
13'b1101100111001,
13'b1101100111010,
13'b1101100111011,
13'b1101100111100,
13'b1101100111101,
13'b1101101001000,
13'b1101101001001,
13'b1101101001010,
13'b1101101001011,
13'b1101101001100,
13'b1101101001101,
13'b1101101011100,
13'b1101101011101,
13'b1110100101000,
13'b1110100101001,
13'b1110100101010,
13'b1110100111000,
13'b1110100111001,
13'b1110100111010,
13'b1110100111011,
13'b1110100111100: edge_mask_reg_512p3[440] <= 1'b1;
 		default: edge_mask_reg_512p3[440] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b11011111000,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100111,
13'b100110101000,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100111,
13'b101110101000,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100111,
13'b111100100100,
13'b111100100101,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000011,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000010,
13'b1010110000011,
13'b1011100100011,
13'b1011100100100,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101100000,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1100101010000,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101100000,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1100101110000,
13'b1100101110001,
13'b1100101110011: edge_mask_reg_512p3[441] <= 1'b1;
 		default: edge_mask_reg_512p3[441] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011111000,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b111100100100,
13'b111100100101,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101000111,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001100110110,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101000110,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1011100100011,
13'b1011100100100,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1100101010001,
13'b1100101010010,
13'b1100101100010: edge_mask_reg_512p3[442] <= 1'b1;
 		default: edge_mask_reg_512p3[442] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011111000,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110110,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b100111001000,
13'b100111001001,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100100,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110100,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111001000,
13'b101111010110,
13'b101111010111,
13'b101111011000,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010011,
13'b110110010100,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100011,
13'b110110100100,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b110110110100,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110110111000,
13'b110110111001,
13'b110111000100,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111001000,
13'b110111010100,
13'b110111010110,
13'b110111010111,
13'b110111011000,
13'b111100100100,
13'b111100100101,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110011000,
13'b111110100011,
13'b111110100100,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b111110101000,
13'b111110110011,
13'b111110110100,
13'b111110110101,
13'b111110110110,
13'b111110110111,
13'b111110111000,
13'b111111000011,
13'b111111000100,
13'b111111000101,
13'b111111000110,
13'b111111000111,
13'b111111001000,
13'b111111010011,
13'b111111010100,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110000,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000000,
13'b1000110000001,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010000,
13'b1000110010001,
13'b1000110010010,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100000,
13'b1000110100001,
13'b1000110100010,
13'b1000110100011,
13'b1000110100100,
13'b1000110100101,
13'b1000110100110,
13'b1000110110000,
13'b1000110110001,
13'b1000110110010,
13'b1000110110011,
13'b1000110110100,
13'b1000110110101,
13'b1000110110110,
13'b1000111000000,
13'b1000111000001,
13'b1000111000010,
13'b1000111000011,
13'b1000111000100,
13'b1000111000101,
13'b1000111010011,
13'b1000111010100,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101110000,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000000,
13'b1001110000001,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010000,
13'b1001110010001,
13'b1001110010010,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1001110100000,
13'b1001110100001,
13'b1001110100010,
13'b1001110100011,
13'b1001110100100,
13'b1001110100101,
13'b1001110110000,
13'b1001110110001,
13'b1001110110010,
13'b1001110110011,
13'b1001110110100,
13'b1001110110101,
13'b1001111000000,
13'b1001111000001,
13'b1001111000010,
13'b1001111000011,
13'b1001111000100,
13'b1001111000101,
13'b1001111010010,
13'b1001111010011,
13'b1001111010100,
13'b1010100100010,
13'b1010100100011,
13'b1010100100100,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010100110101,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100000,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110000,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000000,
13'b1010110000001,
13'b1010110000010,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110010000,
13'b1010110010001,
13'b1010110010010,
13'b1010110010011,
13'b1010110010100,
13'b1010110100000,
13'b1010110100001,
13'b1010110100010,
13'b1010110100011,
13'b1010110100100,
13'b1010110110000,
13'b1010110110001,
13'b1010110110010,
13'b1010110110011,
13'b1010110110100,
13'b1010111000000,
13'b1010111000001,
13'b1010111000010,
13'b1010111000011,
13'b1010111000100,
13'b1010111010010,
13'b1010111010011,
13'b1011100100011,
13'b1011100100100,
13'b1011100110000,
13'b1011100110001,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000000,
13'b1011101000001,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101010000,
13'b1011101010001,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101100000,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101110000,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011110000000,
13'b1011110000001,
13'b1011110000010,
13'b1011110000011,
13'b1011110000100,
13'b1011110010000,
13'b1011110010001,
13'b1011110010010,
13'b1011110010011,
13'b1011110010100,
13'b1011110100000,
13'b1011110100001,
13'b1011110100010,
13'b1011110100011,
13'b1011110100100,
13'b1011110110000,
13'b1011110110001,
13'b1011110110010,
13'b1011110110011,
13'b1011111000000,
13'b1011111000010,
13'b1011111000011: edge_mask_reg_512p3[443] <= 1'b1;
 		default: edge_mask_reg_512p3[443] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110011,
13'b111010110100,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000011,
13'b111011000100,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100011000,
13'b111100011001,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011100011,
13'b1000011100100,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1000011110110,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011101001,
13'b1001011110100,
13'b1001011110110,
13'b1001011110111,
13'b1001011111000,
13'b1001011111001,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100010111,
13'b1001100011000,
13'b1001100011001,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011101001,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010011111000,
13'b1010011111001,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100001001,
13'b1010100010111,
13'b1010100011000,
13'b1010100011001,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100011,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011101000,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011011111000,
13'b1011100000100,
13'b1011100000101,
13'b1011100000110,
13'b1011100000111,
13'b1011100001000,
13'b1011100001001,
13'b1011100010111,
13'b1011100011000,
13'b1011100011001,
13'b1100010100101,
13'b1100010100110,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1100011110111,
13'b1100011111000,
13'b1100100000100,
13'b1100100000101,
13'b1100100000110,
13'b1100100000111,
13'b1100100001000,
13'b1100100010101,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1101011000110,
13'b1101011000111,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1101011100101,
13'b1101011100110,
13'b1101011100111,
13'b1101011101000,
13'b1101011110100,
13'b1101011110101,
13'b1101011110110,
13'b1101011110111,
13'b1101011111000,
13'b1101100000100,
13'b1101100000101,
13'b1101100000110,
13'b1101100000111,
13'b1101100001000,
13'b1101100010101,
13'b1101100010111,
13'b1101100011000,
13'b1110100000101,
13'b1110100000110,
13'b1110100000111,
13'b1110100001000: edge_mask_reg_512p3[444] <= 1'b1;
 		default: edge_mask_reg_512p3[444] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[445] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010101,
13'b110001010110,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000000101,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000000100,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000010100,
13'b1100000010101,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000000100,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1101000010011,
13'b1101000010100,
13'b1101000100010,
13'b1101000100011,
13'b1101000100100,
13'b1110000000000,
13'b1110000000001,
13'b1110000000010,
13'b1110000000011,
13'b1110000000100,
13'b1110000010000,
13'b1110000010001,
13'b1110000010010,
13'b1110000010011,
13'b1110000010100,
13'b1110000100011,
13'b1111000000000,
13'b1111000000001,
13'b1111000000010,
13'b1111000000011,
13'b1111000010000,
13'b1111000010001,
13'b1111000010010: edge_mask_reg_512p3[446] <= 1'b1;
 		default: edge_mask_reg_512p3[446] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110111,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000000110,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1011000000011,
13'b1011000000100,
13'b1011000000101,
13'b1011000000110,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000010110,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1100000000010,
13'b1100000000011,
13'b1100000000100,
13'b1100000000101,
13'b1100000010010,
13'b1100000010011,
13'b1100000010100,
13'b1100000010101,
13'b1100000010110,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000100110,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100000110110,
13'b1100001000100,
13'b1100001000101,
13'b1100001000110,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000000100,
13'b1101000000101,
13'b1101000010010,
13'b1101000010011,
13'b1101000010100,
13'b1101000010101,
13'b1101000100010,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000100110,
13'b1101000110010,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101000110110,
13'b1101001000100,
13'b1101001000101,
13'b1101001000110,
13'b1110000000001,
13'b1110000000010,
13'b1110000000011,
13'b1110000000100,
13'b1110000000101,
13'b1110000010001,
13'b1110000010010,
13'b1110000010011,
13'b1110000010100,
13'b1110000010101,
13'b1110000100001,
13'b1110000100010,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000110010,
13'b1110000110011,
13'b1110000110100,
13'b1110000110101,
13'b1110000110110,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1111000000001,
13'b1111000000010,
13'b1111000000011,
13'b1111000010001,
13'b1111000010010,
13'b1111000010011,
13'b1111000010100,
13'b1111000100001,
13'b1111000100010,
13'b1111000100011,
13'b1111000100100,
13'b1111000110010,
13'b1111000110011,
13'b1111000110100,
13'b1111000110101,
13'b1111001000010,
13'b1111001000011,
13'b1111001000100: edge_mask_reg_512p3[447] <= 1'b1;
 		default: edge_mask_reg_512p3[447] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b1001100100,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110100,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b11001000011,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11010000101,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b101000100001,
13'b101000100010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b110000100000,
13'b110000100001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000000,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b111000010000,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100000,
13'b111000100001,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110000,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111001000000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001010000,
13'b111001010001,
13'b111001010010,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100000,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110000,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000001000000,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001010000,
13'b1000001010001,
13'b1000001010010,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000110000,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001001000000,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001010000,
13'b1001001010001,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001010000,
13'b1010001010001,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000000101,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000000100,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000010100,
13'b1100000010101,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000000100,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1101000010011,
13'b1101000010100,
13'b1101000100000,
13'b1101000100001,
13'b1101000100010,
13'b1101000100011,
13'b1101000100100,
13'b1101000110010,
13'b1110000000000,
13'b1110000000001,
13'b1110000000010,
13'b1110000000011,
13'b1110000000100,
13'b1110000010000,
13'b1110000010001,
13'b1110000010010,
13'b1110000010011,
13'b1110000010100,
13'b1110000100000,
13'b1110000100001,
13'b1110000100011,
13'b1111000000000,
13'b1111000000001,
13'b1111000000010,
13'b1111000000011,
13'b1111000010000,
13'b1111000010001,
13'b1111000010010: edge_mask_reg_512p3[448] <= 1'b1;
 		default: edge_mask_reg_512p3[448] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b10001010100,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100100,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110100,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001010100,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100100,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110100,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000101,
13'b100010000110,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000101,
13'b101010000110,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110101,
13'b110001110110,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010011,
13'b1000001010100,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000010101,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000000101,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000010101,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1100000000010,
13'b1100000000011,
13'b1100000000100,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000010100,
13'b1100000010101,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100000110100,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1100001000011,
13'b1100001000100,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000000100,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1101000010011,
13'b1101000010100,
13'b1101000100000,
13'b1101000100001,
13'b1101000100010,
13'b1101000100011,
13'b1101000100100,
13'b1101000110000,
13'b1101000110001,
13'b1101000110010,
13'b1101000110011,
13'b1101000110100,
13'b1101001000000,
13'b1101001000001,
13'b1101001000010,
13'b1101001000011,
13'b1101001010000,
13'b1101001010001,
13'b1101001010010,
13'b1101001010011,
13'b1110000000000,
13'b1110000000001,
13'b1110000000010,
13'b1110000000011,
13'b1110000000100,
13'b1110000010000,
13'b1110000010001,
13'b1110000010010,
13'b1110000010011,
13'b1110000010100,
13'b1110000100000,
13'b1110000100001,
13'b1110000100010,
13'b1110000100011,
13'b1110000100100,
13'b1110000110000,
13'b1110000110001,
13'b1110000110010,
13'b1110000110011,
13'b1110001000000,
13'b1110001000001,
13'b1110001000010,
13'b1110001000011,
13'b1110001010000,
13'b1111000000001,
13'b1111000000010,
13'b1111000000011,
13'b1111000010000,
13'b1111000010001,
13'b1111000010010,
13'b1111000010011,
13'b1111000100000,
13'b1111000100001,
13'b1111000100010,
13'b1111000110000,
13'b1111000110001,
13'b1111000110010,
13'b1111001000000,
13'b1111001000001,
13'b1111001000010: edge_mask_reg_512p3[449] <= 1'b1;
 		default: edge_mask_reg_512p3[449] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001000,
13'b11001001001,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010011,
13'b1010000010100,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000010011,
13'b1011000010100: edge_mask_reg_512p3[450] <= 1'b1;
 		default: edge_mask_reg_512p3[450] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001001000,
13'b11001001001,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010011,
13'b1010000010100,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000010011,
13'b1011000010100: edge_mask_reg_512p3[451] <= 1'b1;
 		default: edge_mask_reg_512p3[451] <= 1'b0;
 	endcase

    case({x,y,z})
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001001,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110110111,
13'b101110111000,
13'b101110111001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b110110101001,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111101111000,
13'b111101111001,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110001000,
13'b1000101000100,
13'b1000101000101,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110000111,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101010111,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101100111,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001101110111,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110000111,
13'b1010101000011,
13'b1010101000100,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101010110,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101100111,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010101110111,
13'b1010110000011,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110000111,
13'b1011101000011,
13'b1011101000100,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101010110,
13'b1011101100001,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110001,
13'b1011101110010,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011101110111,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110000111,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101010101,
13'b1100101010110,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101100110,
13'b1100101110001,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100101110110,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101010100,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1101101100100,
13'b1101101100101,
13'b1101101100110,
13'b1101101110001,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1101101110101,
13'b1101101110110,
13'b1101110000100,
13'b1101110000101,
13'b1101110000110,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101100001,
13'b1110101100010,
13'b1110101100011,
13'b1110101100100,
13'b1110101100101,
13'b1110101110001,
13'b1110101110010,
13'b1110101110011,
13'b1110101110100,
13'b1110101110101,
13'b1111101100010,
13'b1111101100011,
13'b1111101100100,
13'b1111101100101,
13'b1111101110010,
13'b1111101110011,
13'b1111101110100,
13'b1111101110101: edge_mask_reg_512p3[452] <= 1'b1;
 		default: edge_mask_reg_512p3[452] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[453] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010011000,
13'b1010011001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b100000110011,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001000011,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010011,
13'b100001010100,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100101,
13'b100001100110,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000101011,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010001001,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111001,
13'b110000111010,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001001,
13'b110001001010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001100011,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000110001,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010011,
13'b1000001010100,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000000101,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000110010,
13'b1010000110011,
13'b1011000000011,
13'b1011000000100,
13'b1011000010011,
13'b1011000010100,
13'b1011000100011: edge_mask_reg_512p3[454] <= 1'b1;
 		default: edge_mask_reg_512p3[454] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[455] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10101001,
13'b10101010,
13'b10101011,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101010,
13'b1010101011,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001011100,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011010,
13'b10010011011,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001001100,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001010,
13'b11010001011,
13'b11010011011,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100000111100,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001001100,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101010,
13'b100001101011,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001011000,
13'b101001011001,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000101010,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000011001,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000101001,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000011000,
13'b1000000011001,
13'b1000000100110,
13'b1000000100111,
13'b1000000101000,
13'b1000000101001,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000000111001,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1000001001001,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001011001,
13'b1001000010101,
13'b1001000010110,
13'b1001000010111,
13'b1001000011000,
13'b1001000100110,
13'b1001000100111,
13'b1001000101000,
13'b1001000110110,
13'b1001000110111,
13'b1001000111000,
13'b1001001000110,
13'b1001001000111,
13'b1001001001000,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1010000000101,
13'b1010000000110,
13'b1010000000111,
13'b1010000010101,
13'b1010000010110,
13'b1010000010111,
13'b1010000011000,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000101000,
13'b1010000110110,
13'b1010000110111,
13'b1010000111000,
13'b1010001000110,
13'b1010001000111,
13'b1010001001000,
13'b1010001010111,
13'b1010001011000,
13'b1011000000100,
13'b1011000000101,
13'b1011000000110,
13'b1011000000111,
13'b1011000010101,
13'b1011000010110,
13'b1011000010111,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110110,
13'b1011000110111,
13'b1011000111000,
13'b1011001000110,
13'b1011001000111,
13'b1100000000100,
13'b1100000000101,
13'b1100000000110,
13'b1100000000111,
13'b1100000010101,
13'b1100000010110,
13'b1100000010111,
13'b1100000100101,
13'b1100000100110,
13'b1100000100111,
13'b1100000110101,
13'b1100000110110,
13'b1100000110111,
13'b1100000111000,
13'b1100001000110,
13'b1100001000111,
13'b1101000000101,
13'b1101000000110,
13'b1101000010101,
13'b1101000010110,
13'b1101000010111,
13'b1101000100101,
13'b1101000100110,
13'b1101000100111,
13'b1101000110101,
13'b1101000110110,
13'b1101000110111,
13'b1101001000110,
13'b1101001000111: edge_mask_reg_512p3[456] <= 1'b1;
 		default: edge_mask_reg_512p3[456] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[457] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110111,
13'b11110111000,
13'b100011111000,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110111,
13'b100110111000,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110111,
13'b101110111000,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b111100100111,
13'b111100101000,
13'b111100110111,
13'b111100111000,
13'b111101000111,
13'b111101001000,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101110111,
13'b111101111000,
13'b111110000111,
13'b111110001000,
13'b1000100110110,
13'b1000100110111,
13'b1000100111000,
13'b1000101000110,
13'b1000101000111,
13'b1000101001000,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000111,
13'b1001100110110,
13'b1001100110111,
13'b1001100111000,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000111,
13'b1001110001000,
13'b1010100100111,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1011100100110,
13'b1011100100111,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1100100100111,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1101100100111,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1110100110101,
13'b1110100110110,
13'b1110100110111,
13'b1110101000101,
13'b1110101000110,
13'b1110101000111,
13'b1110101010101,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110110000110,
13'b1110110000111,
13'b1111100110101,
13'b1111100110110,
13'b1111100110111,
13'b1111101000101,
13'b1111101000110,
13'b1111101000111,
13'b1111101010101,
13'b1111101010110,
13'b1111101010111,
13'b1111101100110,
13'b1111101100111,
13'b1111101101000,
13'b1111101110110,
13'b1111101110111,
13'b1111101111000,
13'b1111110000110,
13'b1111110000111: edge_mask_reg_512p3[458] <= 1'b1;
 		default: edge_mask_reg_512p3[458] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110100110,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110110111,
13'b11110111000,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110110111,
13'b100110111000,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110110111,
13'b101110111000,
13'b110011011000,
13'b110011011001,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110010111,
13'b110110011000,
13'b110110011001,
13'b110110100111,
13'b110110101000,
13'b111011101001,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110111,
13'b111101111000,
13'b111110000111,
13'b111110001000,
13'b1000011101010,
13'b1000011111000,
13'b1000011111001,
13'b1000011111010,
13'b1000100001000,
13'b1000100001001,
13'b1000100001010,
13'b1000100011000,
13'b1000100011001,
13'b1000100011010,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100101010,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101000111,
13'b1000101001000,
13'b1000101001001,
13'b1000101010110,
13'b1000101010111,
13'b1000101011000,
13'b1000101011001,
13'b1000101100110,
13'b1000101100111,
13'b1000101101000,
13'b1000101110110,
13'b1000101110111,
13'b1000101111000,
13'b1000110000111,
13'b1001011101010,
13'b1001011111000,
13'b1001011111001,
13'b1001011111010,
13'b1001100001000,
13'b1001100001001,
13'b1001100001010,
13'b1001100011000,
13'b1001100011001,
13'b1001100011010,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100101010,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001100111010,
13'b1001101000110,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101010110,
13'b1001101010111,
13'b1001101011000,
13'b1001101011001,
13'b1001101100110,
13'b1001101100111,
13'b1001101101000,
13'b1001101101001,
13'b1001101110110,
13'b1001101110111,
13'b1001101111000,
13'b1001110000111,
13'b1001110001000,
13'b1010011101010,
13'b1010011111000,
13'b1010011111001,
13'b1010011111010,
13'b1010100001000,
13'b1010100001001,
13'b1010100001010,
13'b1010100011000,
13'b1010100011001,
13'b1010100011010,
13'b1010100011011,
13'b1010100100111,
13'b1010100101000,
13'b1010100101001,
13'b1010100101010,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010100111010,
13'b1010101000110,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101001010,
13'b1010101010110,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101100110,
13'b1010101100111,
13'b1010101101000,
13'b1010101101001,
13'b1010101110110,
13'b1010101110111,
13'b1010101111000,
13'b1010110000110,
13'b1010110000111,
13'b1010110001000,
13'b1011011101001,
13'b1011011101010,
13'b1011011111000,
13'b1011011111001,
13'b1011011111010,
13'b1011100001000,
13'b1011100001001,
13'b1011100001010,
13'b1011100011000,
13'b1011100011001,
13'b1011100011010,
13'b1011100011011,
13'b1011100100111,
13'b1011100101000,
13'b1011100101001,
13'b1011100101010,
13'b1011100110111,
13'b1011100111000,
13'b1011100111001,
13'b1011100111010,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101001001,
13'b1011101001010,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101011001,
13'b1011101100110,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1011101110110,
13'b1011101110111,
13'b1011101111000,
13'b1011110000110,
13'b1011110000111,
13'b1011110001000,
13'b1100011101010,
13'b1100011111001,
13'b1100011111010,
13'b1100011111011,
13'b1100100001000,
13'b1100100001001,
13'b1100100001010,
13'b1100100001011,
13'b1100100011000,
13'b1100100011001,
13'b1100100011010,
13'b1100100011011,
13'b1100100100111,
13'b1100100101000,
13'b1100100101001,
13'b1100100101010,
13'b1100100101011,
13'b1100100110111,
13'b1100100111000,
13'b1100100111001,
13'b1100100111010,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101001001,
13'b1100101001010,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101011001,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101101001,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100110000110,
13'b1100110000111,
13'b1100110001000,
13'b1101011101010,
13'b1101011111001,
13'b1101011111010,
13'b1101011111011,
13'b1101100001000,
13'b1101100001001,
13'b1101100001010,
13'b1101100001011,
13'b1101100011000,
13'b1101100011001,
13'b1101100011010,
13'b1101100011011,
13'b1101100100111,
13'b1101100101000,
13'b1101100101001,
13'b1101100101010,
13'b1101100101011,
13'b1101100110111,
13'b1101100111000,
13'b1101100111001,
13'b1101100111010,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101001001,
13'b1101101001010,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101011001,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101101001,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101110000110,
13'b1101110000111,
13'b1101110001000,
13'b1110011111001,
13'b1110011111010,
13'b1110011111011,
13'b1110100001000,
13'b1110100001001,
13'b1110100001010,
13'b1110100001011,
13'b1110100011000,
13'b1110100011001,
13'b1110100011010,
13'b1110100011011,
13'b1110100100111,
13'b1110100101000,
13'b1110100101001,
13'b1110100101010,
13'b1110100101011,
13'b1110100110111,
13'b1110100111000,
13'b1110100111001,
13'b1110100111010,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101001001,
13'b1110101001010,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101011001,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101101001,
13'b1110101110110,
13'b1110101110111,
13'b1110101111000,
13'b1110110000110,
13'b1110110000111,
13'b1111011111001,
13'b1111011111010,
13'b1111011111011,
13'b1111100001001,
13'b1111100001010,
13'b1111100001011,
13'b1111100011000,
13'b1111100011001,
13'b1111100011010,
13'b1111100011011,
13'b1111100100111,
13'b1111100101000,
13'b1111100101001,
13'b1111100101010,
13'b1111100110111,
13'b1111100111000,
13'b1111100111001,
13'b1111100111010,
13'b1111101000110,
13'b1111101000111,
13'b1111101001000,
13'b1111101001001,
13'b1111101001010,
13'b1111101010110,
13'b1111101010111,
13'b1111101011000,
13'b1111101011001,
13'b1111101100110,
13'b1111101100111,
13'b1111101101000,
13'b1111101101001,
13'b1111101110110,
13'b1111101110111,
13'b1111101111000,
13'b1111110000110,
13'b1111110000111: edge_mask_reg_512p3[459] <= 1'b1;
 		default: edge_mask_reg_512p3[459] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[460] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010111,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010110,
13'b100001010111,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000110,
13'b110001000111,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000100110,
13'b111000100111,
13'b1000000010110,
13'b1000000010111,
13'b1000000011000,
13'b1001000010110,
13'b1001000010111,
13'b1001000011000,
13'b1010000000110,
13'b1010000000111,
13'b1010000001000,
13'b1010000001001,
13'b1010000010110,
13'b1010000010111,
13'b1010000011000,
13'b1010000100110,
13'b1010000100111,
13'b1011000000110,
13'b1011000000111,
13'b1011000001000,
13'b1011000001001,
13'b1011000010110,
13'b1011000010111,
13'b1011000011000,
13'b1011000100110,
13'b1011000100111,
13'b1100000000110,
13'b1100000000111,
13'b1100000001000,
13'b1100000001001,
13'b1100000010110,
13'b1100000010111,
13'b1100000011000,
13'b1100000100111,
13'b1101000000100,
13'b1101000000101,
13'b1101000000110,
13'b1101000000111,
13'b1101000001000,
13'b1101000001001,
13'b1101000001010,
13'b1101000010100,
13'b1101000010101,
13'b1101000010110,
13'b1101000010111,
13'b1101000011000,
13'b1101000100110,
13'b1101000100111,
13'b1110000000100,
13'b1110000000101,
13'b1110000000110,
13'b1110000000111,
13'b1110000001000,
13'b1110000001001,
13'b1110000001010,
13'b1110000010100,
13'b1110000010101,
13'b1110000010110,
13'b1110000010111,
13'b1110000011000,
13'b1110000100110,
13'b1111000000100,
13'b1111000000101,
13'b1111000000110,
13'b1111000000111,
13'b1111000001000,
13'b1111000001001,
13'b1111000010100,
13'b1111000010101,
13'b1111000010110,
13'b1111000010111,
13'b1111000011000,
13'b1111000100110: edge_mask_reg_512p3[461] <= 1'b1;
 		default: edge_mask_reg_512p3[461] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11001000100,
13'b11001000101,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100001000100,
13'b100001000101,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101001000100,
13'b101001000101,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b111000010011,
13'b111000010100,
13'b1000000010010,
13'b1000000010011,
13'b1001000010010,
13'b1001000010011,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010010,
13'b1010000010011,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000000100,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000010001,
13'b1101000010010,
13'b1110000000000,
13'b1110000000001,
13'b1110000000010,
13'b1110000000011,
13'b1111000000000: edge_mask_reg_512p3[462] <= 1'b1;
 		default: edge_mask_reg_512p3[462] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010101,
13'b101010110,
13'b101010111,
13'b101100101,
13'b101100110,
13'b101100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101100101,
13'b1101100110,
13'b1101100111,
13'b1101110101,
13'b1101110110,
13'b1101110111,
13'b1110000101,
13'b1110000110,
13'b1110000111,
13'b1110010101,
13'b1110010110,
13'b1110010111,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110100101,
13'b10110100110,
13'b10110100111,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110110101,
13'b11110110110,
13'b11110110111,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011000,
13'b100110100101,
13'b100110100110,
13'b100110100111,
13'b100110101000,
13'b100110110101,
13'b100110110110,
13'b100110110111,
13'b100111000101,
13'b100111000110,
13'b100111000111,
13'b101100000101,
13'b101100000110,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110100101,
13'b101110100110,
13'b101110100111,
13'b101110101000,
13'b101110110101,
13'b101110110110,
13'b101110110111,
13'b101111000101,
13'b101111000110,
13'b101111000111,
13'b101111010101,
13'b101111010110,
13'b101111010111,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110010101,
13'b110110010110,
13'b110110010111,
13'b110110011000,
13'b110110100101,
13'b110110100110,
13'b110110100111,
13'b110110110101,
13'b110110110110,
13'b110110110111,
13'b110111000101,
13'b110111000110,
13'b110111000111,
13'b110111010110,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010101,
13'b111110010110,
13'b111110010111,
13'b111110100101,
13'b111110100110,
13'b111110100111,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1000110100101,
13'b1000110100110,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001101110110,
13'b1001110000100,
13'b1001110000101,
13'b1001110000110,
13'b1001110010100,
13'b1001110010101,
13'b1001110010110,
13'b1001110100101,
13'b1001110100110,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101000101,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101100110,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010101110110,
13'b1010110000100,
13'b1010110000101,
13'b1010110000110,
13'b1010110010100,
13'b1010110010101,
13'b1010110010110,
13'b1010110100101,
13'b1011100110010,
13'b1011100110011,
13'b1011100110100,
13'b1011101000010,
13'b1011101000011,
13'b1011101000100,
13'b1011101000101,
13'b1011101010010,
13'b1011101010011,
13'b1011101010100,
13'b1011101010101,
13'b1011101100010,
13'b1011101100011,
13'b1011101100100,
13'b1011101100101,
13'b1011101100110,
13'b1011101110011,
13'b1011101110100,
13'b1011101110101,
13'b1011101110110,
13'b1011110000011,
13'b1011110000100,
13'b1011110000101,
13'b1011110000110,
13'b1011110010100,
13'b1011110010101,
13'b1011110010110,
13'b1011110100101,
13'b1011110100110,
13'b1100100110010,
13'b1100100110011,
13'b1100100110100,
13'b1100101000001,
13'b1100101000010,
13'b1100101000011,
13'b1100101000100,
13'b1100101000101,
13'b1100101010001,
13'b1100101010010,
13'b1100101010011,
13'b1100101010100,
13'b1100101010101,
13'b1100101100001,
13'b1100101100010,
13'b1100101100011,
13'b1100101100100,
13'b1100101100101,
13'b1100101110001,
13'b1100101110010,
13'b1100101110011,
13'b1100101110100,
13'b1100101110101,
13'b1100101110110,
13'b1100110000010,
13'b1100110000011,
13'b1100110000100,
13'b1100110000101,
13'b1100110000110,
13'b1100110010100,
13'b1100110010101,
13'b1100110010110,
13'b1100110100100,
13'b1100110100101,
13'b1100110100110,
13'b1101100110010,
13'b1101100110011,
13'b1101101000001,
13'b1101101000010,
13'b1101101000011,
13'b1101101000100,
13'b1101101010000,
13'b1101101010001,
13'b1101101010010,
13'b1101101010011,
13'b1101101010100,
13'b1101101010101,
13'b1101101100000,
13'b1101101100001,
13'b1101101100010,
13'b1101101100011,
13'b1101101100100,
13'b1101101100101,
13'b1101101110001,
13'b1101101110010,
13'b1101101110011,
13'b1101101110100,
13'b1101101110101,
13'b1101110000001,
13'b1101110000010,
13'b1101110000011,
13'b1101110000100,
13'b1101110000101,
13'b1101110000110,
13'b1101110010010,
13'b1101110010011,
13'b1101110010100,
13'b1101110010101,
13'b1101110010110,
13'b1101110100010,
13'b1101110100011,
13'b1101110100100,
13'b1101110100101,
13'b1101110100110,
13'b1110100110010,
13'b1110100110011,
13'b1110101000010,
13'b1110101000011,
13'b1110101000100,
13'b1110101010000,
13'b1110101010001,
13'b1110101010010,
13'b1110101010011,
13'b1110101010100,
13'b1110101100000,
13'b1110101100001,
13'b1110101100010,
13'b1110101100011,
13'b1110101100100,
13'b1110101100101,
13'b1110101110001,
13'b1110101110010,
13'b1110101110011,
13'b1110101110100,
13'b1110101110101,
13'b1110110000001,
13'b1110110000010,
13'b1110110000011,
13'b1110110000100,
13'b1110110000101,
13'b1110110000110,
13'b1110110010010,
13'b1110110010011,
13'b1110110010100,
13'b1110110010101,
13'b1110110010110,
13'b1110110100010,
13'b1110110100011,
13'b1110110100100,
13'b1110110100101,
13'b1110110100110,
13'b1110110110011,
13'b1110110110100,
13'b1111101010001,
13'b1111101010010,
13'b1111101010011,
13'b1111101010100,
13'b1111101100001,
13'b1111101100010,
13'b1111101100011,
13'b1111101100100,
13'b1111101100101,
13'b1111101110001,
13'b1111101110010,
13'b1111101110011,
13'b1111101110100,
13'b1111101110101,
13'b1111110000001,
13'b1111110000010,
13'b1111110000011,
13'b1111110000100,
13'b1111110000101,
13'b1111110000110,
13'b1111110010010,
13'b1111110010011,
13'b1111110010100,
13'b1111110010101,
13'b1111110010110,
13'b1111110100010,
13'b1111110100011,
13'b1111110100100,
13'b1111110100101,
13'b1111110100110,
13'b1111110110011,
13'b1111110110100: edge_mask_reg_512p3[463] <= 1'b1;
 		default: edge_mask_reg_512p3[463] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100111000,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b100001111000,
13'b100001111001,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100111,
13'b100100101000,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100111,
13'b101100101000,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010111,
13'b110100011000,
13'b111010101000,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b1000010101000,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110101,
13'b1000011110110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011101000,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011101000,
13'b1010011110101,
13'b1010011110110,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100011,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011101000,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1100010100111,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000011,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010011,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100011,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1101010100111,
13'b1101010110101,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000011,
13'b1101011000100,
13'b1101011000101,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010011,
13'b1101011010100,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011100101,
13'b1101011100110,
13'b1101011100111,
13'b1101011101000,
13'b1101011110100,
13'b1101011110101,
13'b1101011110110,
13'b1110010110101,
13'b1110010110110,
13'b1110010110111,
13'b1110011000011,
13'b1110011000100,
13'b1110011000101,
13'b1110011000110,
13'b1110011000111,
13'b1110011001000,
13'b1110011010010,
13'b1110011010011,
13'b1110011010100,
13'b1110011010101,
13'b1110011010110,
13'b1110011010111,
13'b1110011011000,
13'b1110011100010,
13'b1110011100011,
13'b1110011100100,
13'b1110011100101,
13'b1110011100110,
13'b1110011100111,
13'b1110011110011,
13'b1110011110100,
13'b1110011110101,
13'b1111010110101,
13'b1111010110110,
13'b1111011000011,
13'b1111011000100,
13'b1111011000101,
13'b1111011000110,
13'b1111011000111,
13'b1111011010010,
13'b1111011010011,
13'b1111011010100,
13'b1111011010101,
13'b1111011010110,
13'b1111011010111,
13'b1111011100010,
13'b1111011100011,
13'b1111011100100,
13'b1111011100101,
13'b1111011110010,
13'b1111011110011: edge_mask_reg_512p3[464] <= 1'b1;
 		default: edge_mask_reg_512p3[464] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b101000101000,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011001,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011101000,
13'b110011101001,
13'b110011111000,
13'b110011111001,
13'b111001010110,
13'b111001010111,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011101000,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010011000,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011100111,
13'b1000011101000,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011100111,
13'b1001011101000,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011100111,
13'b1010011101000,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010000111,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011100111,
13'b1011011101000,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001100010,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1100001110010,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010000110,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010010110,
13'b1100010010111,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010100111,
13'b1100010110101,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000101,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1101001010100,
13'b1101001100010,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001110001,
13'b1101001110010,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101001110110,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1101010000110,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010010101,
13'b1101010010110,
13'b1101010010111,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010100110,
13'b1101010100111,
13'b1101010110100,
13'b1101010110101,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000100,
13'b1101011000101,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1101011100110,
13'b1101011100111,
13'b1110001100010,
13'b1110001100011,
13'b1110001110010,
13'b1110001110011,
13'b1110001110100,
13'b1110001110101,
13'b1110010000010,
13'b1110010000011,
13'b1110010000100,
13'b1110010000101,
13'b1110010000110,
13'b1110010010010,
13'b1110010010011,
13'b1110010010100,
13'b1110010010101,
13'b1110010010110,
13'b1110010100011,
13'b1110010100100,
13'b1110010100101,
13'b1110010100110,
13'b1110010100111,
13'b1110010110011,
13'b1110010110100,
13'b1110010110101,
13'b1110010110110,
13'b1110010110111,
13'b1110011000100,
13'b1110011000101,
13'b1110011000110,
13'b1110011000111,
13'b1110011001000,
13'b1110011010100,
13'b1110011010101,
13'b1110011010110,
13'b1110011010111,
13'b1110011011000,
13'b1110011100110,
13'b1110011100111,
13'b1111001100010,
13'b1111001110010,
13'b1111001110011,
13'b1111010000010,
13'b1111010000011,
13'b1111010000100,
13'b1111010010010,
13'b1111010010011,
13'b1111010010100,
13'b1111010010101,
13'b1111010100011,
13'b1111010100100,
13'b1111010100101,
13'b1111010100110,
13'b1111010110011,
13'b1111010110100,
13'b1111010110101,
13'b1111010110110,
13'b1111011000100,
13'b1111011000101,
13'b1111011000110,
13'b1111011000111,
13'b1111011010100,
13'b1111011010101,
13'b1111011010110,
13'b1111011010111: edge_mask_reg_512p3[465] <= 1'b1;
 		default: edge_mask_reg_512p3[465] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101101000,
13'b101101001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101011001,
13'b10101011010,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101011001,
13'b11101011010,
13'b100001111000,
13'b100001111001,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001001,
13'b100101001010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100111001,
13'b101100111010,
13'b110010011000,
13'b110010011001,
13'b110010101000,
13'b110010101001,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b111010101000,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000111,
13'b111011001000,
13'b111011001001,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011100111,
13'b111011101000,
13'b111011101001,
13'b111011101010,
13'b111011111000,
13'b111011111001,
13'b111011111010,
13'b111100001000,
13'b111100001001,
13'b111100001010,
13'b111100011000,
13'b111100011001,
13'b111100011010,
13'b1000010101000,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1000011101010,
13'b1000011110111,
13'b1000011111000,
13'b1000011111001,
13'b1000011111010,
13'b1000100001000,
13'b1000100001001,
13'b1000100001010,
13'b1000100011000,
13'b1000100011001,
13'b1000100011010,
13'b1001010101000,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011100111,
13'b1001011101000,
13'b1001011101001,
13'b1001011110111,
13'b1001011111000,
13'b1001011111001,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100011000,
13'b1001100011001,
13'b1010010100111,
13'b1010010101000,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1010011100111,
13'b1010011101000,
13'b1010011101001,
13'b1010011110111,
13'b1010011111000,
13'b1010011111001,
13'b1010100000111,
13'b1010100001000,
13'b1010100001001,
13'b1010100010111,
13'b1010100011000,
13'b1010100011001,
13'b1011010100111,
13'b1011010101000,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011010110,
13'b1011011010111,
13'b1011011011000,
13'b1011011011001,
13'b1011011100110,
13'b1011011100111,
13'b1011011101000,
13'b1011011101001,
13'b1011011110111,
13'b1011011111000,
13'b1011011111001,
13'b1011100000111,
13'b1011100001000,
13'b1011100001001,
13'b1011100010111,
13'b1011100011000,
13'b1011100011001,
13'b1100010100111,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100011000110,
13'b1100011000111,
13'b1100011001000,
13'b1100011010110,
13'b1100011010111,
13'b1100011011000,
13'b1100011011001,
13'b1100011100110,
13'b1100011100111,
13'b1100011101000,
13'b1100011101001,
13'b1100011110111,
13'b1100011111000,
13'b1100011111001,
13'b1100100000111,
13'b1100100001000,
13'b1100100001001,
13'b1100100010111,
13'b1100100011000,
13'b1100100011001,
13'b1101010100111,
13'b1101010110110,
13'b1101010110111,
13'b1101010111000,
13'b1101011000101,
13'b1101011000110,
13'b1101011000111,
13'b1101011001000,
13'b1101011010101,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1101011100110,
13'b1101011100111,
13'b1101011101000,
13'b1101011101001,
13'b1101011110110,
13'b1101011110111,
13'b1101011111000,
13'b1101011111001,
13'b1101100000111,
13'b1101100001000,
13'b1101100001001,
13'b1101100010111,
13'b1101100011000,
13'b1101100011001,
13'b1110010110110,
13'b1110010110111,
13'b1110011000100,
13'b1110011000101,
13'b1110011000110,
13'b1110011000111,
13'b1110011001000,
13'b1110011010100,
13'b1110011010101,
13'b1110011010110,
13'b1110011010111,
13'b1110011011000,
13'b1110011100101,
13'b1110011100110,
13'b1110011100111,
13'b1110011101000,
13'b1110011110110,
13'b1110011110111,
13'b1110011111000,
13'b1110100000110,
13'b1110100000111,
13'b1110100001000,
13'b1111010110101,
13'b1111010110110,
13'b1111011000100,
13'b1111011000101,
13'b1111011000110,
13'b1111011000111,
13'b1111011010100,
13'b1111011010101,
13'b1111011010110,
13'b1111011010111,
13'b1111011100101,
13'b1111011100110,
13'b1111011100111,
13'b1111011101000,
13'b1111011110101,
13'b1111011110110,
13'b1111011110111,
13'b1111011111000,
13'b1111100000110,
13'b1111100000111,
13'b1111100001000: edge_mask_reg_512p3[466] <= 1'b1;
 		default: edge_mask_reg_512p3[466] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100110,
13'b10100111,
13'b10110110,
13'b10110111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100110,
13'b1010100111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100110,
13'b100010100111,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010110,
13'b101010010111,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010110,
13'b110010010111,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010101,
13'b1000001010110,
13'b1000001100101,
13'b1000001100110,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100101,
13'b1001001100110,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100101,
13'b1010001100110,
13'b1011000010100,
13'b1011000010101,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1100000010011,
13'b1100000010100,
13'b1100000010101,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100000110110,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001000110,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001100100,
13'b1100001100101,
13'b1100001100110,
13'b1101000010011,
13'b1101000010100,
13'b1101000010101,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000110010,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101001000010,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001000110,
13'b1101001010010,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001010110,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001100110,
13'b1110000010011,
13'b1110000010100,
13'b1110000010101,
13'b1110000100010,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000110010,
13'b1110000110011,
13'b1110000110100,
13'b1110000110101,
13'b1110001000010,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1110001000110,
13'b1110001010010,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001010110,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001100110,
13'b1111000100010,
13'b1111000100011,
13'b1111000100100,
13'b1111000100101,
13'b1111000110010,
13'b1111000110011,
13'b1111000110100,
13'b1111000110101,
13'b1111001000010,
13'b1111001000011,
13'b1111001000100,
13'b1111001000101,
13'b1111001010010,
13'b1111001010011,
13'b1111001010100,
13'b1111001010101,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001100101,
13'b1111001100110: edge_mask_reg_512p3[467] <= 1'b1;
 		default: edge_mask_reg_512p3[467] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100110,
13'b10100111,
13'b10110110,
13'b10110111,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100110,
13'b1010100111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100110,
13'b100010100111,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010110,
13'b101010010111,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010110,
13'b110010010111,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000010111,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100101,
13'b1001001100110,
13'b1010000000100,
13'b1010000000101,
13'b1010000000110,
13'b1010000000111,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000010111,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100101,
13'b1010001100110,
13'b1011000000100,
13'b1011000000101,
13'b1011000000110,
13'b1011000000111,
13'b1011000010100,
13'b1011000010101,
13'b1011000010110,
13'b1011000010111,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1100000000100,
13'b1100000000101,
13'b1100000000110,
13'b1100000010100,
13'b1100000010101,
13'b1100000010110,
13'b1100000100100,
13'b1100000100101,
13'b1100000100110,
13'b1100000110100,
13'b1100000110101,
13'b1100000110110,
13'b1100001000100,
13'b1100001000101,
13'b1100001000110,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001100100,
13'b1100001100101,
13'b1100001100110,
13'b1101000000010,
13'b1101000000011,
13'b1101000000100,
13'b1101000000101,
13'b1101000000110,
13'b1101000010010,
13'b1101000010011,
13'b1101000010100,
13'b1101000010101,
13'b1101000010110,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000100110,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101000110110,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001000110,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001010110,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001100110,
13'b1110000000010,
13'b1110000000011,
13'b1110000000100,
13'b1110000000101,
13'b1110000000110,
13'b1110000010010,
13'b1110000010011,
13'b1110000010100,
13'b1110000010101,
13'b1110000010110,
13'b1110000100010,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000100110,
13'b1110000110010,
13'b1110000110011,
13'b1110000110100,
13'b1110000110101,
13'b1110000110110,
13'b1110001000010,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1110001000110,
13'b1110001010010,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001010110,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001100110,
13'b1111000000010,
13'b1111000000011,
13'b1111000000100,
13'b1111000000101,
13'b1111000000110,
13'b1111000010010,
13'b1111000010011,
13'b1111000010100,
13'b1111000010101,
13'b1111000010110,
13'b1111000100010,
13'b1111000100011,
13'b1111000100100,
13'b1111000100101,
13'b1111000100110,
13'b1111000110010,
13'b1111000110011,
13'b1111000110100,
13'b1111000110101,
13'b1111000110110,
13'b1111001000010,
13'b1111001000011,
13'b1111001000100,
13'b1111001000101,
13'b1111001000110,
13'b1111001010010,
13'b1111001010011,
13'b1111001010100,
13'b1111001010101,
13'b1111001010110,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001100101,
13'b1111001100110: edge_mask_reg_512p3[468] <= 1'b1;
 		default: edge_mask_reg_512p3[468] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100110,
13'b10100111,
13'b10110110,
13'b10110111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100110,
13'b1010100111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010100110,
13'b100010100111,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010110,
13'b101010010111,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010110,
13'b110010010111,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100101,
13'b1000001100110,
13'b1001000010011,
13'b1001000010100,
13'b1001000010101,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1011000010010,
13'b1011000010011,
13'b1011000010100,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1100000010010,
13'b1100000010011,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000100100,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001100100,
13'b1100001100101,
13'b1100001100110,
13'b1101000010010,
13'b1101000010011,
13'b1101000100001,
13'b1101000100010,
13'b1101000100011,
13'b1101000100100,
13'b1101000110000,
13'b1101000110001,
13'b1101000110010,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101001000000,
13'b1101001000001,
13'b1101001000010,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001010000,
13'b1101001010001,
13'b1101001010010,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001010110,
13'b1101001100001,
13'b1101001100010,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001100110,
13'b1110000100011,
13'b1110000110000,
13'b1110000110001,
13'b1110000110010,
13'b1110000110011,
13'b1110000110100,
13'b1110000110101,
13'b1110001000000,
13'b1110001000001,
13'b1110001000010,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1110001010001,
13'b1110001010010,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001010110,
13'b1110001100001,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001100110,
13'b1111000110100,
13'b1111001000001,
13'b1111001000010,
13'b1111001000011,
13'b1111001000100,
13'b1111001000101,
13'b1111001010001,
13'b1111001010010,
13'b1111001010011,
13'b1111001010100,
13'b1111001010101,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001100101,
13'b1111001100110: edge_mask_reg_512p3[469] <= 1'b1;
 		default: edge_mask_reg_512p3[469] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110110,
13'b11011110111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110110,
13'b100011110111,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110110,
13'b101011110111,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100110,
13'b110011100111,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b1000000110101,
13'b1000000110110,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000100,
13'b1000011000101,
13'b1001000110101,
13'b1001000110110,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000100,
13'b1001011000101,
13'b1010000110101,
13'b1010000110110,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000100,
13'b1010011000101,
13'b1011000110100,
13'b1011000110101,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1100000110100,
13'b1100000110101,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1100001100110,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010000110,
13'b1100010010001,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010100001,
13'b1100010100010,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010110001,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100010110101,
13'b1100011000011,
13'b1100011000100,
13'b1101000110100,
13'b1101000110101,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001010010,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001010110,
13'b1101001100010,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001100110,
13'b1101001110001,
13'b1101001110010,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101001110110,
13'b1101010000001,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1101010010001,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010010101,
13'b1101010100001,
13'b1101010100010,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010110001,
13'b1101010110010,
13'b1101010110011,
13'b1101010110100,
13'b1101010110101,
13'b1101011000011,
13'b1101011000100,
13'b1110000110100,
13'b1110000110101,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1110001010010,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001010110,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001100110,
13'b1110001110001,
13'b1110001110010,
13'b1110001110011,
13'b1110001110100,
13'b1110001110101,
13'b1110001110110,
13'b1110010000001,
13'b1110010000010,
13'b1110010000011,
13'b1110010000100,
13'b1110010000101,
13'b1110010010001,
13'b1110010010010,
13'b1110010010011,
13'b1110010010100,
13'b1110010010101,
13'b1110010100001,
13'b1110010100010,
13'b1110010100011,
13'b1110010100100,
13'b1110010100101,
13'b1110010110001,
13'b1110010110010,
13'b1110010110011,
13'b1110010110100,
13'b1110010110101,
13'b1110011000011,
13'b1110011000100,
13'b1111001000011,
13'b1111001000100,
13'b1111001000101,
13'b1111001010010,
13'b1111001010011,
13'b1111001010100,
13'b1111001010101,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001100101,
13'b1111001100110,
13'b1111001110001,
13'b1111001110010,
13'b1111001110011,
13'b1111001110100,
13'b1111001110101,
13'b1111010000001,
13'b1111010000010,
13'b1111010000011,
13'b1111010000100,
13'b1111010000101,
13'b1111010010001,
13'b1111010010010,
13'b1111010010011,
13'b1111010010100,
13'b1111010010101,
13'b1111010100001,
13'b1111010100010,
13'b1111010100011,
13'b1111010110001,
13'b1111010110010: edge_mask_reg_512p3[470] <= 1'b1;
 		default: edge_mask_reg_512p3[470] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100111,
13'b11011101000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100111,
13'b100011101000,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100111,
13'b101011101000,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010111,
13'b110011011000,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110111,
13'b111010111000,
13'b1000000110101,
13'b1000000110110,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000010000110,
13'b1000010000111,
13'b1000010001000,
13'b1000010001001,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010111000,
13'b1001000110101,
13'b1001000110110,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010001001,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010111000,
13'b1010000110101,
13'b1010000110110,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001010111,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001101000,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010001001,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010111000,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001010111,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001100111,
13'b1011001101000,
13'b1011001110101,
13'b1011001110110,
13'b1011001110111,
13'b1011001111000,
13'b1011010000110,
13'b1011010000111,
13'b1011010001000,
13'b1011010001001,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010011001,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010111000,
13'b1011010111001,
13'b1100000110100,
13'b1100000110101,
13'b1100001000100,
13'b1100001000101,
13'b1100001000110,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001010111,
13'b1100001100100,
13'b1100001100101,
13'b1100001100110,
13'b1100001100111,
13'b1100001101000,
13'b1100001110101,
13'b1100001110110,
13'b1100001110111,
13'b1100001111000,
13'b1100010000101,
13'b1100010000110,
13'b1100010000111,
13'b1100010001000,
13'b1100010001001,
13'b1100010010110,
13'b1100010010111,
13'b1100010011000,
13'b1100010011001,
13'b1100010100111,
13'b1100010101000,
13'b1100010101001,
13'b1100010111000,
13'b1100010111001,
13'b1101000110100,
13'b1101000110101,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001000110,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001010110,
13'b1101001010111,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001100110,
13'b1101001100111,
13'b1101001101000,
13'b1101001110100,
13'b1101001110101,
13'b1101001110110,
13'b1101001110111,
13'b1101001111000,
13'b1101010000101,
13'b1101010000110,
13'b1101010000111,
13'b1101010001000,
13'b1101010001001,
13'b1101010010110,
13'b1101010010111,
13'b1101010011000,
13'b1101010011001,
13'b1101010011010,
13'b1101010100111,
13'b1101010101000,
13'b1101010101001,
13'b1101010101010,
13'b1101010111000,
13'b1101010111001,
13'b1110000110100,
13'b1110000110101,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1110001000110,
13'b1110001010010,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001010110,
13'b1110001010111,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001100110,
13'b1110001100111,
13'b1110001101000,
13'b1110001110010,
13'b1110001110011,
13'b1110001110100,
13'b1110001110101,
13'b1110001110110,
13'b1110001110111,
13'b1110001111000,
13'b1110010000100,
13'b1110010000101,
13'b1110010000110,
13'b1110010000111,
13'b1110010001000,
13'b1110010001001,
13'b1110010010110,
13'b1110010010111,
13'b1110010011000,
13'b1110010011001,
13'b1110010011010,
13'b1110010100111,
13'b1110010101000,
13'b1110010101001,
13'b1110010101010,
13'b1110010111000,
13'b1110010111001,
13'b1111001000011,
13'b1111001000100,
13'b1111001000101,
13'b1111001000110,
13'b1111001010010,
13'b1111001010011,
13'b1111001010100,
13'b1111001010101,
13'b1111001010110,
13'b1111001010111,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001100101,
13'b1111001100110,
13'b1111001100111,
13'b1111001110010,
13'b1111001110011,
13'b1111001110100,
13'b1111001110101,
13'b1111001110110,
13'b1111001110111,
13'b1111001111000,
13'b1111010000011,
13'b1111010000100,
13'b1111010000101,
13'b1111010000110,
13'b1111010000111,
13'b1111010001000,
13'b1111010001001,
13'b1111010010101,
13'b1111010010110,
13'b1111010010111,
13'b1111010011000,
13'b1111010011001,
13'b1111010100110,
13'b1111010100111,
13'b1111010101000,
13'b1111010101001,
13'b1111010111000,
13'b1111010111001: edge_mask_reg_512p3[471] <= 1'b1;
 		default: edge_mask_reg_512p3[471] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10100111,
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010011,
13'b11010100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100011,
13'b11100100,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110001,
13'b11110010,
13'b11110011,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000001,
13'b100000010,
13'b100000011,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010001,
13'b100010010,
13'b100010011,
13'b100010100,
13'b100010101,
13'b100010111,
13'b100011000,
13'b100100001,
13'b100100010,
13'b100100011,
13'b100100100,
13'b100100111,
13'b100101000,
13'b100110001,
13'b100110010,
13'b100110011,
13'b100110100,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000001,
13'b101000010,
13'b101000011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010001,
13'b101010010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010011,
13'b1011010100,
13'b1011010101,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100011,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110001,
13'b1011110010,
13'b1011110011,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000001,
13'b1100000010,
13'b1100000011,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010001,
13'b1100010010,
13'b1100010011,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100001,
13'b1100100010,
13'b1100100011,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110001,
13'b1100110010,
13'b1100110011,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000001,
13'b1101000010,
13'b1101000011,
13'b1101000100,
13'b1101000101,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010001,
13'b1101010010,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010111,
13'b10011011000,
13'b10011011010,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010001,
13'b10100010010,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100001,
13'b10100100010,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110001,
13'b10100110010,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000001,
13'b10101000010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010011,
13'b11011010100,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010011,
13'b11101010100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010: edge_mask_reg_512p3[472] <= 1'b1;
 		default: edge_mask_reg_512p3[472] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10101000,
13'b10101001,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010011,
13'b11010100,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100011,
13'b11100100,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110001,
13'b11110010,
13'b11110011,
13'b11110100,
13'b11110101,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000001,
13'b100000010,
13'b100000011,
13'b100000100,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100010001,
13'b100010010,
13'b100010011,
13'b100010100,
13'b100010101,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100001,
13'b100100010,
13'b100100011,
13'b100100100,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110001,
13'b100110010,
13'b100110011,
13'b100110100,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000001,
13'b101000010,
13'b101000011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010001,
13'b101010010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100001,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010011,
13'b1011010100,
13'b1011010101,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100011,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110001,
13'b1011110010,
13'b1011110011,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000001,
13'b1100000010,
13'b1100000011,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010001,
13'b1100010010,
13'b1100010011,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100100001,
13'b1100100010,
13'b1100100011,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100110001,
13'b1100110010,
13'b1100110011,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000001,
13'b1101000010,
13'b1101000011,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010001,
13'b1101010010,
13'b1101010011,
13'b1101010100,
13'b1101010101,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100001,
13'b1101100010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010001,
13'b10100010010,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100001,
13'b10100100010,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110001,
13'b10100110010,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000001,
13'b10101000010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010001,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100001,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110001,
13'b10101110010,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100001,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110001,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000001,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010001,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100001,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110001,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000011,
13'b100100000100,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110001,
13'b100100110010,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000001,
13'b100101000010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010001,
13'b100101010010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100001,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110001,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000001,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110111001,
13'b100110111010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110011,
13'b101100110100,
13'b101100110110,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101010001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110001,
13'b101101110010,
13'b101101110011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000001,
13'b101110000010,
13'b101110000011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010011,
13'b101110010100,
13'b101110010101,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111001,
13'b101110111010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010011,
13'b110101010100,
13'b110101011001,
13'b110101011010,
13'b110101100001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101101001,
13'b110101101010,
13'b110101110001,
13'b110101110010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101111001,
13'b110101111010,
13'b110110000011,
13'b110110000100,
13'b110110000101,
13'b110110000110: edge_mask_reg_512p3[473] <= 1'b1;
 		default: edge_mask_reg_512p3[473] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110110,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101011000,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b100001101001,
13'b100001101010,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101010111011,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011001011,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b110010001001,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010010,
13'b111011010011,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111011111001,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010101000,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000011110111,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100000111,
13'b1000100010010,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100000110,
13'b1001100000111,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100010110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010011110101,
13'b1010011110110,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100000100,
13'b1010100000101,
13'b1010100000110,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100010100,
13'b1010100010101,
13'b1010100010110,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1011100000100,
13'b1011100000101,
13'b1011100010011,
13'b1011100010100,
13'b1011100010101,
13'b1100010100101,
13'b1100010100110,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011010011,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011100011,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1100011110011,
13'b1100011110100,
13'b1100011110101,
13'b1100100000011,
13'b1100100000100,
13'b1100100000101,
13'b1100100010011,
13'b1100100010100,
13'b1100100010101: edge_mask_reg_512p3[474] <= 1'b1;
 		default: edge_mask_reg_512p3[474] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110101,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100000,
13'b10010100001,
13'b10010100010,
13'b10010100011,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110010,
13'b10010110011,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000000,
13'b11010000001,
13'b11010000010,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010000,
13'b11010010001,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100000,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110000,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000000,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000000,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010000,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100000,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110000,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000000,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110110,
13'b100100110111,
13'b101001100101,
13'b101001100110,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000000,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110110,
13'b101100110111,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010000,
13'b110010010001,
13'b110010010010,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010000,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100100110,
13'b110100100111,
13'b111010100000,
13'b111010100001,
13'b111010100010,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000000,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010000,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b1000010110000,
13'b1000010110001,
13'b1000010110010,
13'b1000011000000,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011010000,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010011,
13'b1001010110000,
13'b1001011000000,
13'b1001011000001,
13'b1001011000010,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100010010,
13'b1010011000000,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100010010,
13'b1011011000000,
13'b1011011010000,
13'b1011011010001,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011100000001,
13'b1011100000010,
13'b1011100000011,
13'b1100011010000,
13'b1100011100000,
13'b1100011100001,
13'b1100011110000,
13'b1100011110001,
13'b1101011100000: edge_mask_reg_512p3[475] <= 1'b1;
 		default: edge_mask_reg_512p3[475] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11110101,
13'b11110110,
13'b11110111,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b101000101,
13'b101000110,
13'b101000111,
13'b101010110,
13'b101010111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101010110,
13'b1101010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010000,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010100000,
13'b10010100001,
13'b10010100010,
13'b10010100011,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010110010,
13'b10010110011,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000000,
13'b11010000001,
13'b11010000010,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010000,
13'b11010010001,
13'b11010010010,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100000,
13'b11010100001,
13'b11010100010,
13'b11010100011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110000,
13'b11010110001,
13'b11010110010,
13'b11010110011,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000000,
13'b11011000001,
13'b11011000010,
13'b11011000011,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010010,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100010000000,
13'b100010000001,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010000,
13'b100010010001,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100000,
13'b100010100001,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110000,
13'b100010110001,
13'b100010110010,
13'b100010110011,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000000,
13'b100011000001,
13'b100011000010,
13'b100011000011,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010000,
13'b100011010001,
13'b100011010010,
13'b100011010011,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100000,
13'b100011100001,
13'b100011100010,
13'b100011100011,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110010,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b101001100101,
13'b101001100110,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101010000000,
13'b101010000001,
13'b101010000010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010000,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100000,
13'b101010100001,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110000,
13'b101010110001,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000000,
13'b101011000001,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010000,
13'b101011010001,
13'b101011010010,
13'b101011010011,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100000,
13'b101011100001,
13'b101011100010,
13'b101011100011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110000,
13'b101011110001,
13'b101011110010,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101100000001,
13'b101100000010,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101101000110,
13'b101101000111,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010010000,
13'b110010010001,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010100000,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010110000,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110011000000,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010000,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011100000,
13'b110011100001,
13'b110011100010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110000,
13'b110011110001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110101000110,
13'b110101000111,
13'b111010100000,
13'b111010100001,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110000,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000000,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010000,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010110,
13'b111011010111,
13'b111011100000,
13'b111011100001,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b1000010110000,
13'b1000010110001,
13'b1000011000000,
13'b1000011000001,
13'b1000011000010,
13'b1000011010000,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100100011,
13'b1001011000000,
13'b1001011010000,
13'b1001011010001,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100100001,
13'b1001100100010,
13'b1010011010000,
13'b1010011100000,
13'b1010011100001,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100010001,
13'b1010100010010,
13'b1011011100000,
13'b1011011110000,
13'b1011100000000: edge_mask_reg_512p3[476] <= 1'b1;
 		default: edge_mask_reg_512p3[476] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[477] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101101100,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001001,
13'b101110001010,
13'b101110001011,
13'b101110011010,
13'b101110101010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001001,
13'b110110001010,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110001001,
13'b111110001010,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101011010,
13'b1000101101000,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1000110001001,
13'b1000110001010,
13'b1000110001011,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100011001,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001100111010,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101001010,
13'b1001101011000,
13'b1001101011001,
13'b1001101011010,
13'b1001101101000,
13'b1001101101001,
13'b1001101101010,
13'b1001101111001,
13'b1001101111010,
13'b1001101111011,
13'b1001110001001,
13'b1001110001010,
13'b1001110001011,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1010100011001,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100101001,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101001010,
13'b1010101011000,
13'b1010101011001,
13'b1010101011010,
13'b1010101101000,
13'b1010101101001,
13'b1010101101010,
13'b1010101111001,
13'b1010101111010,
13'b1010101111011,
13'b1010110001001,
13'b1010110001010,
13'b1010110001011,
13'b1011100000110,
13'b1011100000111,
13'b1011100001000,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100101001,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011100111001,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101001001,
13'b1011101001010,
13'b1011101010111,
13'b1011101011000,
13'b1011101011001,
13'b1011101011010,
13'b1011101101000,
13'b1011101101001,
13'b1011101101010,
13'b1011101111000,
13'b1011101111001,
13'b1011101111010,
13'b1011101111011,
13'b1011110001001,
13'b1011110001010,
13'b1100100000110,
13'b1100100000111,
13'b1100100001000,
13'b1100100010101,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100101001,
13'b1100100110100,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100100111001,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101001001,
13'b1100101001010,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101011001,
13'b1100101011010,
13'b1100101100111,
13'b1100101101000,
13'b1100101101001,
13'b1100101101010,
13'b1100101101011,
13'b1100101111000,
13'b1100101111001,
13'b1100101111010,
13'b1100101111011,
13'b1100110001001,
13'b1100110001010,
13'b1100110001011,
13'b1101100010101,
13'b1101100010110,
13'b1101100010111,
13'b1101100011000,
13'b1101100100100,
13'b1101100100101,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101100111001,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101001001,
13'b1101101001010,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101011001,
13'b1101101011010,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101101001,
13'b1101101101010,
13'b1101101110111,
13'b1101101111000,
13'b1101101111001,
13'b1101101111010,
13'b1101110001000,
13'b1101110001001,
13'b1101110001010,
13'b1110100100100,
13'b1110100100101,
13'b1110100100110,
13'b1110100110101,
13'b1110100110110,
13'b1110100110111,
13'b1110100111000,
13'b1110101000101,
13'b1110101000110,
13'b1110101000111,
13'b1110101001000,
13'b1110101001001,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101011001,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101101001,
13'b1110101101010,
13'b1110101110111,
13'b1110101111000,
13'b1110101111001,
13'b1110101111010,
13'b1110110000111,
13'b1110110001000,
13'b1110110001001,
13'b1111100110101,
13'b1111100110110,
13'b1111101000101,
13'b1111101000110,
13'b1111101000111,
13'b1111101010110,
13'b1111101010111,
13'b1111101011000,
13'b1111101100110,
13'b1111101100111,
13'b1111101101000,
13'b1111101101001,
13'b1111101110111,
13'b1111101111000,
13'b1111101111001,
13'b1111110000111,
13'b1111110001000: edge_mask_reg_512p3[478] <= 1'b1;
 		default: edge_mask_reg_512p3[478] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b10110101100,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110101100,
13'b11110111010,
13'b11110111011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100100111100,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101001100,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101011100,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110011010,
13'b100110011011,
13'b100110101010,
13'b100110101011,
13'b101011101001,
13'b101011101010,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101100111011,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101001011,
13'b101101011001,
13'b101101011010,
13'b101101011011,
13'b101101101001,
13'b101101101010,
13'b101101101011,
13'b101101111001,
13'b101101111010,
13'b101101111011,
13'b101110001010,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101011011,
13'b110101101001,
13'b110101101010,
13'b110101101011,
13'b110101111001,
13'b110101111010,
13'b110101111011,
13'b110110001010,
13'b111100000111,
13'b111100001000,
13'b111100001001,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100101010,
13'b111100111000,
13'b111100111001,
13'b111100111010,
13'b111101001000,
13'b111101001001,
13'b111101001010,
13'b111101011000,
13'b111101011001,
13'b111101011010,
13'b111101011011,
13'b111101101001,
13'b111101101010,
13'b111101101011,
13'b111101111001,
13'b111101111010,
13'b111101111011,
13'b111110001001,
13'b111110001010,
13'b1000100000111,
13'b1000100001000,
13'b1000100001001,
13'b1000100010111,
13'b1000100011000,
13'b1000100011001,
13'b1000100100111,
13'b1000100101000,
13'b1000100101001,
13'b1000100110111,
13'b1000100111000,
13'b1000100111001,
13'b1000100111010,
13'b1000101001000,
13'b1000101001001,
13'b1000101001010,
13'b1000101011000,
13'b1000101011001,
13'b1000101011010,
13'b1000101101001,
13'b1000101101010,
13'b1000101101011,
13'b1000101111001,
13'b1000101111010,
13'b1000101111011,
13'b1000110001001,
13'b1000110001010,
13'b1001100000110,
13'b1001100000111,
13'b1001100001000,
13'b1001100001001,
13'b1001100010110,
13'b1001100010111,
13'b1001100011000,
13'b1001100011001,
13'b1001100100111,
13'b1001100101000,
13'b1001100101001,
13'b1001100110111,
13'b1001100111000,
13'b1001100111001,
13'b1001100111010,
13'b1001101000111,
13'b1001101001000,
13'b1001101001001,
13'b1001101001010,
13'b1001101011000,
13'b1001101011001,
13'b1001101011010,
13'b1001101101000,
13'b1001101101001,
13'b1001101101010,
13'b1001101101011,
13'b1001101111001,
13'b1001101111010,
13'b1001101111011,
13'b1001110001001,
13'b1001110001010,
13'b1010100000110,
13'b1010100000111,
13'b1010100001000,
13'b1010100010110,
13'b1010100010111,
13'b1010100011000,
13'b1010100011001,
13'b1010100100110,
13'b1010100100111,
13'b1010100101000,
13'b1010100101001,
13'b1010100110110,
13'b1010100110111,
13'b1010100111000,
13'b1010100111001,
13'b1010100111010,
13'b1010101000111,
13'b1010101001000,
13'b1010101001001,
13'b1010101001010,
13'b1010101010111,
13'b1010101011000,
13'b1010101011001,
13'b1010101011010,
13'b1010101101000,
13'b1010101101001,
13'b1010101101010,
13'b1010101111000,
13'b1010101111001,
13'b1010101111010,
13'b1010110001001,
13'b1011100000110,
13'b1011100000111,
13'b1011100001000,
13'b1011100010101,
13'b1011100010110,
13'b1011100010111,
13'b1011100011000,
13'b1011100100100,
13'b1011100100101,
13'b1011100100110,
13'b1011100100111,
13'b1011100101000,
13'b1011100101001,
13'b1011100110101,
13'b1011100110110,
13'b1011100110111,
13'b1011100111000,
13'b1011100111001,
13'b1011101000110,
13'b1011101000111,
13'b1011101001000,
13'b1011101001001,
13'b1011101001010,
13'b1011101010110,
13'b1011101010111,
13'b1011101011000,
13'b1011101011001,
13'b1011101011010,
13'b1011101100111,
13'b1011101101000,
13'b1011101101001,
13'b1011101101010,
13'b1011101110111,
13'b1011101111000,
13'b1011101111001,
13'b1011101111010,
13'b1011110001001,
13'b1100100000110,
13'b1100100000111,
13'b1100100001000,
13'b1100100010101,
13'b1100100010110,
13'b1100100010111,
13'b1100100011000,
13'b1100100100100,
13'b1100100100101,
13'b1100100100110,
13'b1100100100111,
13'b1100100101000,
13'b1100100101001,
13'b1100100110100,
13'b1100100110101,
13'b1100100110110,
13'b1100100110111,
13'b1100100111000,
13'b1100100111001,
13'b1100101000101,
13'b1100101000110,
13'b1100101000111,
13'b1100101001000,
13'b1100101001001,
13'b1100101001010,
13'b1100101010101,
13'b1100101010110,
13'b1100101010111,
13'b1100101011000,
13'b1100101011001,
13'b1100101011010,
13'b1100101100110,
13'b1100101100111,
13'b1100101101000,
13'b1100101101001,
13'b1100101101010,
13'b1100101110110,
13'b1100101110111,
13'b1100101111000,
13'b1100101111001,
13'b1100101111010,
13'b1100110000111,
13'b1101100010101,
13'b1101100010110,
13'b1101100010111,
13'b1101100011000,
13'b1101100100100,
13'b1101100100101,
13'b1101100100110,
13'b1101100100111,
13'b1101100101000,
13'b1101100110101,
13'b1101100110110,
13'b1101100110111,
13'b1101100111000,
13'b1101100111001,
13'b1101101000101,
13'b1101101000110,
13'b1101101000111,
13'b1101101001000,
13'b1101101001001,
13'b1101101010101,
13'b1101101010110,
13'b1101101010111,
13'b1101101011000,
13'b1101101011001,
13'b1101101011010,
13'b1101101100110,
13'b1101101100111,
13'b1101101101000,
13'b1101101101001,
13'b1101101101010,
13'b1101101110110,
13'b1101101110111,
13'b1101101111000,
13'b1101101111001,
13'b1101101111010,
13'b1101110000111,
13'b1110100100100,
13'b1110100100101,
13'b1110100100110,
13'b1110100110101,
13'b1110100110110,
13'b1110100110111,
13'b1110101000101,
13'b1110101000110,
13'b1110101000111,
13'b1110101010110,
13'b1110101010111,
13'b1110101011000,
13'b1110101100110,
13'b1110101100111,
13'b1110101101000,
13'b1110101110111,
13'b1110101111000: edge_mask_reg_512p3[479] <= 1'b1;
 		default: edge_mask_reg_512p3[479] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000111,
13'b1100001000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b100001010111,
13'b100001011000,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b101001010111,
13'b101001011000,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111010111001,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010011,
13'b1001010000010,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010010001,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010100000,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010110000,
13'b1010010110001,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010010001,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010100000,
13'b1011010100001,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010110000,
13'b1011010110001,
13'b1011010110010,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1100010000011,
13'b1100010000100,
13'b1100010010001,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010100001,
13'b1100010100010,
13'b1100010100011,
13'b1100010100100,
13'b1100010110001,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100011000011,
13'b1100011000100,
13'b1101010010001,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010100001,
13'b1101010100010,
13'b1101010100011,
13'b1101010100100,
13'b1101010110001,
13'b1101010110010,
13'b1101010110011,
13'b1101010110100,
13'b1110010010001,
13'b1110010010010,
13'b1110010010011,
13'b1110010100001,
13'b1110010100010,
13'b1110010100011,
13'b1110010110001,
13'b1110010110010,
13'b1110010110011,
13'b1111010010010,
13'b1111010100010,
13'b1111010110010: edge_mask_reg_512p3[480] <= 1'b1;
 		default: edge_mask_reg_512p3[480] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100110000110,
13'b100110000111,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101110000110,
13'b101110000111,
13'b110011100111,
13'b110011101000,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1010100000010,
13'b1010100000011,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101010001,
13'b1010101010010: edge_mask_reg_512p3[481] <= 1'b1;
 		default: edge_mask_reg_512p3[481] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101100110,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100011000,
13'b1100101000,
13'b1100110111,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110111,
13'b11101111000,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110111,
13'b100101111000,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100010000,
13'b101100010001,
13'b101100010010,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000000,
13'b110100000001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100111,
13'b110101101000,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100011001,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100101001,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1001100000000,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000010,
13'b1001101000011,
13'b1010100000010,
13'b1010100000011,
13'b1010100010000,
13'b1010100010010,
13'b1010100010011,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011: edge_mask_reg_512p3[482] <= 1'b1;
 		default: edge_mask_reg_512p3[482] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100110110,
13'b100110111,
13'b100111000,
13'b100111001,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110010110,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110100111,
13'b11110101000,
13'b11110101001,
13'b11110101010,
13'b11110110111,
13'b11110111000,
13'b11110111001,
13'b11110111010,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110010111,
13'b100110011000,
13'b100110011001,
13'b100110011010,
13'b100110100111,
13'b100110101000,
13'b100110101001,
13'b100110101010,
13'b100110110111,
13'b100110111000,
13'b100110111001,
13'b100110111010,
13'b100111001000,
13'b100111001001,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110010101,
13'b101110010110,
13'b101110010111,
13'b101110011000,
13'b101110011001,
13'b101110011010,
13'b101110100111,
13'b101110101000,
13'b101110101001,
13'b101110101010,
13'b101110111000,
13'b101110111001,
13'b110011100111,
13'b110011101000,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101101010,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b110101111010,
13'b110110000100,
13'b110110000101,
13'b110110000110,
13'b110110000111,
13'b110110001000,
13'b110110001001,
13'b110110001010,
13'b110110010101,
13'b110110010110,
13'b110110011000,
13'b110110011001,
13'b110110101000,
13'b110110101001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101001000,
13'b111101001001,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101010111,
13'b111101011000,
13'b111101011001,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101100111,
13'b111101101000,
13'b111101101001,
13'b111101110010,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b111101110110,
13'b111101110111,
13'b111110000011,
13'b111110000100,
13'b111110000101,
13'b111110000110,
13'b111110000111,
13'b111110010011,
13'b111110010100,
13'b111110010101,
13'b111110010110,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010000,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101010111,
13'b1000101100000,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101100110,
13'b1000101100111,
13'b1000101110001,
13'b1000101110010,
13'b1000101110011,
13'b1000101110100,
13'b1000101110101,
13'b1000101110110,
13'b1000110000010,
13'b1000110000011,
13'b1000110000100,
13'b1000110000101,
13'b1000110000110,
13'b1000110010011,
13'b1000110010100,
13'b1000110010101,
13'b1000110010110,
13'b1001100000000,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000000,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101000101,
13'b1001101010000,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101010101,
13'b1001101010110,
13'b1001101100000,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1001101100101,
13'b1001101100110,
13'b1001101110001,
13'b1001101110010,
13'b1001101110011,
13'b1001101110100,
13'b1001101110101,
13'b1001110000010,
13'b1001110000011,
13'b1001110000100,
13'b1001110000101,
13'b1001110010011,
13'b1001110010100,
13'b1001110010101,
13'b1010100000010,
13'b1010100000011,
13'b1010100010000,
13'b1010100010010,
13'b1010100010011,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100110000,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010100110100,
13'b1010101000000,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101000100,
13'b1010101010000,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1010101010100,
13'b1010101010101,
13'b1010101100001,
13'b1010101100010,
13'b1010101100011,
13'b1010101100100,
13'b1010101100101,
13'b1010101110001,
13'b1010101110010,
13'b1010101110011,
13'b1010101110100,
13'b1010101110101,
13'b1010110000011,
13'b1010110000100: edge_mask_reg_512p3[483] <= 1'b1;
 		default: edge_mask_reg_512p3[483] <= 1'b0;
 	endcase

    case({x,y,z})
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b1110000110,
13'b1110000111,
13'b1110001000,
13'b1110010111,
13'b1110011000,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100110000,
13'b100100110001,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100110000111,
13'b100110001000,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010000,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100000,
13'b101100100001,
13'b101100100010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110000,
13'b101100110001,
13'b101100110010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000000,
13'b101101000001,
13'b101101000010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100010,
13'b101101100011,
13'b101101100100,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101110000111,
13'b101110001000,
13'b110011100111,
13'b110011101000,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010000,
13'b110100010001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100000,
13'b110100100001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110000,
13'b110100110001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000000,
13'b110101000001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101010001,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101100010,
13'b110101100011,
13'b110101100100,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110111,
13'b110101111000,
13'b110101111001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111100111001,
13'b111101000000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101001000,
13'b111101001001,
13'b111101010001,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101100010,
13'b111101100011,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000000,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101010010,
13'b1000101010011,
13'b1000101100010,
13'b1000101100011,
13'b1001100000000,
13'b1001100000010,
13'b1001100000011,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000010,
13'b1001101000011,
13'b1010100000010,
13'b1010100000011,
13'b1010100010000,
13'b1010100010010,
13'b1010100010011,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011: edge_mask_reg_512p3[484] <= 1'b1;
 		default: edge_mask_reg_512p3[484] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b101010110,
13'b101010111,
13'b101011000,
13'b101100110,
13'b101100111,
13'b101101000,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101100110,
13'b1101100111,
13'b1101101000,
13'b1101110110,
13'b1101110111,
13'b1101111000,
13'b10010010111,
13'b10010011000,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101110111,
13'b11101111000,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101110111,
13'b100101111000,
13'b101010100111,
13'b101010101000,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000101,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100100010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101010111,
13'b110101011000,
13'b110101100111,
13'b110101101000,
13'b111011000100,
13'b111011000101,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110000,
13'b111011110001,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000000,
13'b111100000001,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100001000,
13'b111100010000,
13'b111100010001,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100011000,
13'b111100100000,
13'b111100100001,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100101000,
13'b111100110000,
13'b111100110001,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111100111000,
13'b111101000001,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b1000011000100,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100000,
13'b1000011100001,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1000011110000,
13'b1000011110001,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000000,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100010000,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100100000,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100110000,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011010000,
13'b1001011010001,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100000,
13'b1001011100001,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110000,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000000,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100010000,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100100000,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100110000,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001101000010,
13'b1001101000011,
13'b1010011000010,
13'b1010011010000,
13'b1010011010001,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011100000,
13'b1010011100001,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011110000,
13'b1010011110001,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1010100000000,
13'b1010100000001,
13'b1010100000010,
13'b1010100000011,
13'b1010100010000,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100100000,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1011011010000,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011100000,
13'b1011011100001,
13'b1011011100010,
13'b1011011100011,
13'b1011011110000,
13'b1011011110001,
13'b1011011110010,
13'b1011011110011,
13'b1011100000000,
13'b1011100000001: edge_mask_reg_512p3[485] <= 1'b1;
 		default: edge_mask_reg_512p3[485] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[486] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011001000,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000101001,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010111000,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000011000,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010110,
13'b111010010111,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010101,
13'b1000010010110,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000010111,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000100111,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010101,
13'b1001010010110,
13'b1010000000101,
13'b1010000000110,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000010111,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000100111,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001010111,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1011000000100,
13'b1011000000101,
13'b1011000000110,
13'b1011000010100,
13'b1011000010101,
13'b1011000010110,
13'b1011000010111,
13'b1011000100011,
13'b1011000100100,
13'b1011000100101,
13'b1011000100110,
13'b1011000100111,
13'b1011000110011,
13'b1011000110100,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001000111,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001010111,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001100111,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011001110111,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1100000000100,
13'b1100000000101,
13'b1100000000110,
13'b1100000010100,
13'b1100000010101,
13'b1100000010110,
13'b1100000100011,
13'b1100000100100,
13'b1100000100101,
13'b1100000100110,
13'b1100000110011,
13'b1100000110100,
13'b1100000110101,
13'b1100000110110,
13'b1100001000011,
13'b1100001000100,
13'b1100001000101,
13'b1100001000110,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1100001100110,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010100,
13'b1101000000100,
13'b1101000000101,
13'b1101000000110,
13'b1101000010100,
13'b1101000010101,
13'b1101000010110,
13'b1101000100011,
13'b1101000100100,
13'b1101000100101,
13'b1101000100110,
13'b1101000110011,
13'b1101000110100,
13'b1101000110101,
13'b1101000110110,
13'b1101001000011,
13'b1101001000100,
13'b1101001000101,
13'b1101001000110,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001010110,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001100110,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101001110110,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1110000000100,
13'b1110000000101,
13'b1110000000110,
13'b1110000010011,
13'b1110000010100,
13'b1110000010101,
13'b1110000010110,
13'b1110000100011,
13'b1110000100100,
13'b1110000100101,
13'b1110000100110,
13'b1110000110011,
13'b1110000110100,
13'b1110000110101,
13'b1110000110110,
13'b1110001000011,
13'b1110001000100,
13'b1110001000101,
13'b1110001000110,
13'b1110001010011,
13'b1110001010100,
13'b1110001010101,
13'b1110001010110,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001100110,
13'b1110001110011,
13'b1110001110100,
13'b1110001110101,
13'b1110010000011,
13'b1110010000100,
13'b1110010000101,
13'b1111000010011,
13'b1111000010100,
13'b1111000010101,
13'b1111000100011,
13'b1111000100100,
13'b1111000100101,
13'b1111000110011,
13'b1111000110100,
13'b1111000110101,
13'b1111001000011,
13'b1111001000100,
13'b1111001000101,
13'b1111001010011,
13'b1111001010100,
13'b1111001010101,
13'b1111001100011,
13'b1111001100100,
13'b1111001100101,
13'b1111001110011,
13'b1111001110100,
13'b1111001110101,
13'b1111010000011,
13'b1111010000100,
13'b1111010000101: edge_mask_reg_512p3[487] <= 1'b1;
 		default: edge_mask_reg_512p3[487] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000111,
13'b11011001000,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011001000,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010110,
13'b111010010111,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010101,
13'b1000010010110,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010010101,
13'b1001010010110,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001110010,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001110010,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011001110111,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010010100,
13'b1011010010101,
13'b1100001010011,
13'b1100001010100,
13'b1100001010101,
13'b1100001100010,
13'b1100001100011,
13'b1100001100100,
13'b1100001100101,
13'b1100001100110,
13'b1100001110010,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010011,
13'b1100010010100,
13'b1101001010011,
13'b1101001010100,
13'b1101001010101,
13'b1101001100010,
13'b1101001100011,
13'b1101001100100,
13'b1101001100101,
13'b1101001100110,
13'b1101001110010,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101001110110,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1110001010011,
13'b1110001010100,
13'b1110001100010,
13'b1110001100011,
13'b1110001100100,
13'b1110001100101,
13'b1110001110010,
13'b1110001110011,
13'b1110001110100,
13'b1110001110101,
13'b1110010000011,
13'b1110010000100,
13'b1110010000101,
13'b1111001100010,
13'b1111001100011,
13'b1111001100100,
13'b1111001110010,
13'b1111001110011,
13'b1111001110100,
13'b1111010000010,
13'b1111010000011,
13'b1111010000100,
13'b1111010000101: edge_mask_reg_512p3[488] <= 1'b1;
 		default: edge_mask_reg_512p3[488] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101100111,
13'b101101000,
13'b101101001,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110010111,
13'b1110011000,
13'b1110011001,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110101000,
13'b11110101001,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110011000,
13'b100110011001,
13'b101010101001,
13'b101010101010,
13'b101010110101,
13'b101010111001,
13'b101010111010,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011011011,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011101011,
13'b101011110011,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100000011,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100010011,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100100011,
13'b101100100100,
13'b101100100101,
13'b101100100110,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100110011,
13'b101100110100,
13'b101100110101,
13'b101100110110,
13'b101100110111,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101000011,
13'b101101000100,
13'b101101000101,
13'b101101000110,
13'b101101000111,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101010011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101010111,
13'b101101011000,
13'b101101011001,
13'b101101011010,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101100111,
13'b101101101000,
13'b101101101001,
13'b101101101010,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111000,
13'b101101111001,
13'b101101111010,
13'b101110000111,
13'b101110001000,
13'b101110001001,
13'b101110001010,
13'b101110011000,
13'b101110011001,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011010,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011110011,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110011111010,
13'b110100000011,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100001010,
13'b110100010011,
13'b110100010100,
13'b110100010101,
13'b110100010110,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100011010,
13'b110100100011,
13'b110100100100,
13'b110100100101,
13'b110100100110,
13'b110100100111,
13'b110100101000,
13'b110100101001,
13'b110100101010,
13'b110100110010,
13'b110100110011,
13'b110100110100,
13'b110100110101,
13'b110100110110,
13'b110100110111,
13'b110100111000,
13'b110100111001,
13'b110100111010,
13'b110101000010,
13'b110101000011,
13'b110101000100,
13'b110101000101,
13'b110101000110,
13'b110101000111,
13'b110101001000,
13'b110101001001,
13'b110101001010,
13'b110101010010,
13'b110101010011,
13'b110101010100,
13'b110101010101,
13'b110101010110,
13'b110101010111,
13'b110101011000,
13'b110101011001,
13'b110101011010,
13'b110101100011,
13'b110101100100,
13'b110101100101,
13'b110101100110,
13'b110101100111,
13'b110101101000,
13'b110101101001,
13'b110101110011,
13'b110101110100,
13'b110101110101,
13'b110101110110,
13'b110101111000,
13'b110101111001,
13'b110110001000,
13'b110110001001,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011100010,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011100111,
13'b111011110010,
13'b111011110011,
13'b111011110100,
13'b111011110101,
13'b111011110110,
13'b111011110111,
13'b111100000010,
13'b111100000011,
13'b111100000100,
13'b111100000101,
13'b111100000110,
13'b111100000111,
13'b111100010010,
13'b111100010011,
13'b111100010100,
13'b111100010101,
13'b111100010110,
13'b111100010111,
13'b111100100010,
13'b111100100011,
13'b111100100100,
13'b111100100101,
13'b111100100110,
13'b111100100111,
13'b111100110010,
13'b111100110011,
13'b111100110100,
13'b111100110101,
13'b111100110110,
13'b111100110111,
13'b111101000010,
13'b111101000011,
13'b111101000100,
13'b111101000101,
13'b111101000110,
13'b111101000111,
13'b111101010010,
13'b111101010011,
13'b111101010100,
13'b111101010101,
13'b111101010110,
13'b111101100010,
13'b111101100011,
13'b111101100100,
13'b111101100101,
13'b111101100110,
13'b111101110011,
13'b111101110100,
13'b111101110101,
13'b1000011000100,
13'b1000011000101,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100010,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110010,
13'b1000011110011,
13'b1000011110100,
13'b1000011110101,
13'b1000011110110,
13'b1000100000001,
13'b1000100000010,
13'b1000100000011,
13'b1000100000100,
13'b1000100000101,
13'b1000100000110,
13'b1000100010001,
13'b1000100010010,
13'b1000100010011,
13'b1000100010100,
13'b1000100010101,
13'b1000100010110,
13'b1000100100001,
13'b1000100100010,
13'b1000100100011,
13'b1000100100100,
13'b1000100100101,
13'b1000100100110,
13'b1000100110001,
13'b1000100110010,
13'b1000100110011,
13'b1000100110100,
13'b1000100110101,
13'b1000100110110,
13'b1000101000001,
13'b1000101000010,
13'b1000101000011,
13'b1000101000100,
13'b1000101000101,
13'b1000101000110,
13'b1000101010001,
13'b1000101010010,
13'b1000101010011,
13'b1000101010100,
13'b1000101010101,
13'b1000101010110,
13'b1000101100001,
13'b1000101100010,
13'b1000101100011,
13'b1000101100100,
13'b1000101100101,
13'b1000101110011,
13'b1000101110100,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011100010,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110001,
13'b1001011110010,
13'b1001011110011,
13'b1001011110100,
13'b1001011110101,
13'b1001100000001,
13'b1001100000010,
13'b1001100000011,
13'b1001100000100,
13'b1001100000101,
13'b1001100010001,
13'b1001100010010,
13'b1001100010011,
13'b1001100010100,
13'b1001100010101,
13'b1001100100001,
13'b1001100100010,
13'b1001100100011,
13'b1001100100100,
13'b1001100100101,
13'b1001100110001,
13'b1001100110010,
13'b1001100110011,
13'b1001100110100,
13'b1001100110101,
13'b1001101000001,
13'b1001101000010,
13'b1001101000011,
13'b1001101000100,
13'b1001101010001,
13'b1001101010010,
13'b1001101010011,
13'b1001101010100,
13'b1001101100001,
13'b1001101100010,
13'b1001101100011,
13'b1001101100100,
13'b1010011010010,
13'b1010011010011,
13'b1010011100010,
13'b1010011100011,
13'b1010011110010,
13'b1010011110011,
13'b1010100000010,
13'b1010100000011,
13'b1010100010001,
13'b1010100010010,
13'b1010100010011,
13'b1010100100001,
13'b1010100100010,
13'b1010100100011,
13'b1010100110001,
13'b1010100110010,
13'b1010100110011,
13'b1010101000001,
13'b1010101000010,
13'b1010101000011,
13'b1010101010001,
13'b1010101010010,
13'b1010101010011,
13'b1011100100010,
13'b1011100110010,
13'b1011101000001,
13'b1011101000010,
13'b1011101010001,
13'b1011101010010: edge_mask_reg_512p3[489] <= 1'b1;
 		default: edge_mask_reg_512p3[489] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[490] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011001,
13'b10011010,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110010,
13'b11110011,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000010,
13'b100000011,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010010,
13'b100010011,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100100010,
13'b100100011,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100110010,
13'b100110011,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b100111100,
13'b101000010,
13'b101000011,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101001100,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101011100,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b101101100,
13'b1010101001,
13'b1010101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010100,
13'b1011010101,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011110010,
13'b1011110011,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100000010,
13'b1100000011,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100010010,
13'b1100010011,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100100010,
13'b1100100011,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100110010,
13'b1100110011,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101000010,
13'b1101000011,
13'b1101000100,
13'b1101000101,
13'b1101000110,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101001100,
13'b1101010010,
13'b1101010011,
13'b1101010100,
13'b1101010101,
13'b1101010110,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101011100,
13'b1101100010,
13'b1101100011,
13'b1101100100,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b1101101100,
13'b1101110010,
13'b1101110011,
13'b1101110111,
13'b1101111000,
13'b1101111001,
13'b1101111010,
13'b1101111011,
13'b1101111100,
13'b1110000010,
13'b1110000011,
13'b1110000111,
13'b1110001000,
13'b1110001001,
13'b1110001010,
13'b1110001011,
13'b1110001100,
13'b1110010010,
13'b1110011000,
13'b1110011001,
13'b1110011010,
13'b1110011011,
13'b1110011100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010010,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100100010,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100110010,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101000010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101001100,
13'b10101010010,
13'b10101010011,
13'b10101010100,
13'b10101010101,
13'b10101010110,
13'b10101010111,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101011100,
13'b10101100010,
13'b10101100011,
13'b10101100100,
13'b10101100101,
13'b10101100110,
13'b10101100111,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101101100,
13'b10101110010,
13'b10101110011,
13'b10101110100,
13'b10101110101,
13'b10101110110,
13'b10101110111,
13'b10101111000,
13'b10101111001,
13'b10101111010,
13'b10101111011,
13'b10101111100,
13'b10110000010,
13'b10110000011,
13'b10110000100,
13'b10110000101,
13'b10110000110,
13'b10110000111,
13'b10110001000,
13'b10110001001,
13'b10110001010,
13'b10110001011,
13'b10110001100,
13'b10110010010,
13'b10110010011,
13'b10110010100,
13'b10110010101,
13'b10110010110,
13'b10110010111,
13'b10110011000,
13'b10110011001,
13'b10110011010,
13'b10110011011,
13'b10110011100,
13'b10110100110,
13'b10110100111,
13'b10110101000,
13'b10110101001,
13'b10110101010,
13'b10110101011,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101000010,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101001100,
13'b11101010010,
13'b11101010011,
13'b11101010100,
13'b11101010101,
13'b11101010110,
13'b11101010111,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101011100,
13'b11101100010,
13'b11101100011,
13'b11101100100,
13'b11101100101,
13'b11101100110,
13'b11101100111,
13'b11101101000,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b11101101100,
13'b11101110010,
13'b11101110011,
13'b11101110100,
13'b11101110101,
13'b11101110110,
13'b11101110111,
13'b11101111000,
13'b11101111001,
13'b11101111010,
13'b11101111011,
13'b11101111100,
13'b11110000010,
13'b11110000011,
13'b11110000100,
13'b11110000101,
13'b11110000110,
13'b11110000111,
13'b11110001000,
13'b11110001001,
13'b11110001010,
13'b11110001011,
13'b11110001100,
13'b11110010010,
13'b11110010011,
13'b11110010100,
13'b11110010101,
13'b11110010110,
13'b11110010111,
13'b11110011000,
13'b11110011001,
13'b11110011010,
13'b11110011011,
13'b11110011100,
13'b11110100100,
13'b11110100101,
13'b11110100110,
13'b11110100111,
13'b11110101001,
13'b11110101010,
13'b11110101011,
13'b11110111001,
13'b11110111010,
13'b11110111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110100,
13'b100011110101,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101000110,
13'b100101000111,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101010011,
13'b100101010100,
13'b100101010101,
13'b100101010110,
13'b100101010111,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101100010,
13'b100101100011,
13'b100101100100,
13'b100101100101,
13'b100101100110,
13'b100101100111,
13'b100101101000,
13'b100101101001,
13'b100101101010,
13'b100101101011,
13'b100101110010,
13'b100101110011,
13'b100101110100,
13'b100101110101,
13'b100101110110,
13'b100101110111,
13'b100101111000,
13'b100101111001,
13'b100101111010,
13'b100101111011,
13'b100110000010,
13'b100110000011,
13'b100110000100,
13'b100110000101,
13'b100110000110,
13'b100110000111,
13'b100110001000,
13'b100110001001,
13'b100110001010,
13'b100110001011,
13'b100110010100,
13'b100110010101,
13'b100110010110,
13'b100110010111,
13'b100110011001,
13'b100110011010,
13'b100110011011,
13'b100110100100,
13'b100110100101,
13'b100110101001,
13'b100110101010,
13'b100110101011,
13'b100110111001,
13'b100110111010,
13'b100110111011,
13'b101011111010,
13'b101011111011,
13'b101100001010,
13'b101100001011,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111010,
13'b101100111011,
13'b101101000100,
13'b101101000101,
13'b101101001010,
13'b101101001011,
13'b101101010100,
13'b101101010101,
13'b101101010110,
13'b101101011010,
13'b101101011011,
13'b101101100100,
13'b101101100101,
13'b101101100110,
13'b101101101010,
13'b101101101011,
13'b101101110100,
13'b101101110101,
13'b101101110110,
13'b101101110111,
13'b101101111010,
13'b101101111011,
13'b101110000100,
13'b101110000101,
13'b101110000110,
13'b101110000111,
13'b101110001010,
13'b101110010100,
13'b101110010101,
13'b101110010110: edge_mask_reg_512p3[491] <= 1'b1;
 		default: edge_mask_reg_512p3[491] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11110001,
13'b11110010,
13'b11110011,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b11111100,
13'b100000001,
13'b100000010,
13'b100000011,
13'b100000100,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100001100,
13'b100010001,
13'b100010010,
13'b100010011,
13'b100010100,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100011100,
13'b100100001,
13'b100100010,
13'b100100011,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100101010,
13'b100101011,
13'b100101100,
13'b100110001,
13'b100110010,
13'b100110011,
13'b100110111,
13'b100111000,
13'b100111001,
13'b100111010,
13'b100111011,
13'b101000001,
13'b101000010,
13'b101000011,
13'b101000111,
13'b101001000,
13'b101001001,
13'b101001010,
13'b101001011,
13'b101010111,
13'b101011000,
13'b101011001,
13'b101011010,
13'b101011011,
13'b101100111,
13'b101101000,
13'b101101001,
13'b101101010,
13'b101101011,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010011,
13'b1011010100,
13'b1011010101,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100011,
13'b1011100100,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011110001,
13'b1011110010,
13'b1011110011,
13'b1011110100,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100000001,
13'b1100000010,
13'b1100000011,
13'b1100000100,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100010001,
13'b1100010010,
13'b1100010011,
13'b1100010100,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100011100,
13'b1100100001,
13'b1100100010,
13'b1100100011,
13'b1100100100,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100101010,
13'b1100101011,
13'b1100101100,
13'b1100110001,
13'b1100110010,
13'b1100110011,
13'b1100110100,
13'b1100110101,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b1100111001,
13'b1100111010,
13'b1100111011,
13'b1100111100,
13'b1101000001,
13'b1101000010,
13'b1101000011,
13'b1101000111,
13'b1101001000,
13'b1101001001,
13'b1101001010,
13'b1101001011,
13'b1101010111,
13'b1101011000,
13'b1101011001,
13'b1101011010,
13'b1101011011,
13'b1101100111,
13'b1101101000,
13'b1101101001,
13'b1101101010,
13'b1101101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011010011,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100011,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011110010,
13'b10011110011,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100000001,
13'b10100000010,
13'b10100000011,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100010001,
13'b10100010010,
13'b10100010011,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100011011,
13'b10100011100,
13'b10100100001,
13'b10100100010,
13'b10100100011,
13'b10100100100,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100101010,
13'b10100101011,
13'b10100101100,
13'b10100110001,
13'b10100110010,
13'b10100110011,
13'b10100110100,
13'b10100110101,
13'b10100110110,
13'b10100110111,
13'b10100111000,
13'b10100111001,
13'b10100111010,
13'b10100111011,
13'b10100111100,
13'b10101000001,
13'b10101000010,
13'b10101000011,
13'b10101000100,
13'b10101000101,
13'b10101000110,
13'b10101000111,
13'b10101001000,
13'b10101001001,
13'b10101001010,
13'b10101001011,
13'b10101010011,
13'b10101010100,
13'b10101011000,
13'b10101011001,
13'b10101011010,
13'b10101011011,
13'b10101101000,
13'b10101101001,
13'b10101101010,
13'b10101101011,
13'b10101111010,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010011,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100011,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110010,
13'b11011110011,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100000010,
13'b11100000011,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100001100,
13'b11100010001,
13'b11100010010,
13'b11100010011,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100011011,
13'b11100011100,
13'b11100100010,
13'b11100100011,
13'b11100100100,
13'b11100100101,
13'b11100100110,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100101010,
13'b11100101011,
13'b11100101100,
13'b11100110010,
13'b11100110011,
13'b11100110100,
13'b11100110101,
13'b11100110110,
13'b11100110111,
13'b11100111000,
13'b11100111001,
13'b11100111010,
13'b11100111011,
13'b11100111100,
13'b11101000011,
13'b11101000100,
13'b11101000101,
13'b11101000110,
13'b11101000111,
13'b11101001000,
13'b11101001001,
13'b11101001010,
13'b11101001011,
13'b11101010011,
13'b11101010100,
13'b11101011000,
13'b11101011001,
13'b11101011010,
13'b11101011011,
13'b11101101001,
13'b11101101010,
13'b11101101011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100100,
13'b100011100101,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011101011,
13'b100011110011,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100011111011,
13'b100011111100,
13'b100100000011,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100001011,
13'b100100001100,
13'b100100010011,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100011011,
13'b100100011100,
13'b100100100011,
13'b100100100100,
13'b100100100101,
13'b100100100110,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100101010,
13'b100100101011,
13'b100100101100,
13'b100100110011,
13'b100100110100,
13'b100100110101,
13'b100100110110,
13'b100100110111,
13'b100100111000,
13'b100100111001,
13'b100100111010,
13'b100100111011,
13'b100101000011,
13'b100101000100,
13'b100101000101,
13'b100101001000,
13'b100101001001,
13'b100101001010,
13'b100101001011,
13'b100101011000,
13'b100101011001,
13'b100101011010,
13'b100101011011,
13'b100101101001,
13'b100101101010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101011111011,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100001011,
13'b101100011000,
13'b101100011001,
13'b101100011010,
13'b101100011011,
13'b101100100100,
13'b101100100101,
13'b101100101000,
13'b101100101001,
13'b101100101010,
13'b101100101011,
13'b101100110100,
13'b101100110101,
13'b101100111000,
13'b101100111001,
13'b101100111010,
13'b101101001000,
13'b101101001001,
13'b101101001010,
13'b101101011001,
13'b101101011010,
13'b110100001001,
13'b110100001010,
13'b110100011001,
13'b110100011010,
13'b110100101001,
13'b110100101010: edge_mask_reg_512p3[492] <= 1'b1;
 		default: edge_mask_reg_512p3[492] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10011100,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10101100,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b10111011,
13'b10111100,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11001011,
13'b11001100,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11011011,
13'b11011100,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11101011,
13'b11101100,
13'b11111000,
13'b11111001,
13'b11111010,
13'b11111011,
13'b100001000,
13'b100001001,
13'b100001010,
13'b100001011,
13'b100011000,
13'b100011001,
13'b100011010,
13'b100011011,
13'b100101001,
13'b100101010,
13'b100101011,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010101100,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1010111100,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011001100,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011011100,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011101011,
13'b1011101100,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1011111011,
13'b1011111100,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100001011,
13'b1100001100,
13'b1100011001,
13'b1100011010,
13'b1100011011,
13'b1100101010,
13'b1100101011,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10010111100,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011001100,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011011100,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011101100,
13'b10011111001,
13'b10011111010,
13'b10011111011,
13'b10011111100,
13'b10100001001,
13'b10100001010,
13'b10100001011,
13'b10100001100,
13'b10100011010,
13'b10100011011,
13'b10100101010,
13'b10100101011,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001011100,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001101100,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11001111100,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010001100,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010011100,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010101100,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11010111100,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011001100,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011011100,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011101100,
13'b11011111001,
13'b11011111010,
13'b11011111011,
13'b11011111100,
13'b11100001001,
13'b11100001010,
13'b11100001011,
13'b11100011010,
13'b11100011011,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010001100,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010011100,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010101100,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100010111100,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011001100,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101010,
13'b100011101011,
13'b100011111010,
13'b100011111011,
13'b101000101001,
13'b101000101010,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101000111011,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001001011,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011001,
13'b101011011010,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110111,
13'b111001111000,
13'b111001111001,
13'b111010000111,
13'b111010001000,
13'b111010001001,
13'b111010001010,
13'b111010010111,
13'b111010011000,
13'b111010011001,
13'b111010011010,
13'b111010100111,
13'b111010101000,
13'b111010101001,
13'b111010101010,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b1000000110111,
13'b1000000111000,
13'b1000000111001,
13'b1000001000111,
13'b1000001001000,
13'b1000001001001,
13'b1000001010111,
13'b1000001011000,
13'b1000001011001,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001101001,
13'b1000001110111,
13'b1000001111000,
13'b1000001111001,
13'b1000010000111,
13'b1000010001000,
13'b1000010001001,
13'b1000010010111,
13'b1000010011000,
13'b1000010011001,
13'b1000010100101,
13'b1000010100111,
13'b1000010101000,
13'b1000010101001,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011011000,
13'b1000011011001,
13'b1000011011010,
13'b1001000110110,
13'b1001000110111,
13'b1001000111000,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001001000,
13'b1001001001001,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1001001011001,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001101001,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001001111001,
13'b1001010000101,
13'b1001010000110,
13'b1001010000111,
13'b1001010001000,
13'b1001010001001,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010011000,
13'b1001010011001,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010101000,
13'b1001010101001,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001010111000,
13'b1001010111001,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010000111000,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001001000,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001101000,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010001111000,
13'b1010001111001,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010000111,
13'b1010010001000,
13'b1010010001001,
13'b1010010010101,
13'b1010010010110,
13'b1010010010111,
13'b1010010011000,
13'b1010010011001,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010101000,
13'b1010010101001,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010010111000,
13'b1010010111001,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1011000110110,
13'b1011000110111,
13'b1011000111000,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001000111,
13'b1011001001000,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001010111,
13'b1011001011000,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001100111,
13'b1011001101000,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011001110111,
13'b1011001111000,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010000111,
13'b1011010001000,
13'b1011010010101,
13'b1011010010110,
13'b1011010010111,
13'b1011010011000,
13'b1011010011001,
13'b1011010100101,
13'b1011010100110,
13'b1011010100111,
13'b1011010101000,
13'b1011010101001,
13'b1011010110101,
13'b1011010110110,
13'b1011010110111,
13'b1011010111000,
13'b1011010111001,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011001000,
13'b1011011001001,
13'b1011011010111,
13'b1011011011000,
13'b1011011011001,
13'b1100000110110,
13'b1100000110111,
13'b1100001000100,
13'b1100001000101,
13'b1100001000110,
13'b1100001000111,
13'b1100001001000,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001010111,
13'b1100001011000,
13'b1100001100100,
13'b1100001100101,
13'b1100001100110,
13'b1100001100111,
13'b1100001101000,
13'b1100001110100,
13'b1100001110101,
13'b1100001110110,
13'b1100001110111,
13'b1100001111000,
13'b1100010000101,
13'b1100010000110,
13'b1100010000111,
13'b1100010001000,
13'b1100010010101,
13'b1100010010110,
13'b1100010010111,
13'b1100010011000,
13'b1100010100110,
13'b1100010100111,
13'b1100010101000,
13'b1100010110110,
13'b1100010110111,
13'b1100010111000,
13'b1100010111001,
13'b1100011000111,
13'b1100011001000,
13'b1100011001001,
13'b1100011011000,
13'b1100011011001: edge_mask_reg_512p3[493] <= 1'b1;
 		default: edge_mask_reg_512p3[493] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11001000,
13'b11001001,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101000111011,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001001011,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101001,
13'b101010101010,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111000111001,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001001001,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001011000,
13'b111001011001,
13'b111001100011,
13'b111001100100,
13'b111001100110,
13'b111001100111,
13'b111001101000,
13'b111001101001,
13'b111001110011,
13'b111001110110,
13'b111001110111,
13'b111001111000,
13'b111010000110,
13'b111010000111,
13'b1000000110110,
13'b1000000110111,
13'b1000000111000,
13'b1000000111001,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001001000,
13'b1000001001001,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001011000,
13'b1000001011001,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001100111,
13'b1000001101000,
13'b1000001101001,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000001110111,
13'b1000001111000,
13'b1000010000110,
13'b1001000110101,
13'b1001000110110,
13'b1001000110111,
13'b1001000111000,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001000111,
13'b1001001001000,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001010111,
13'b1001001011000,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001100110,
13'b1001001100111,
13'b1001001101000,
13'b1001001110011,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001001110111,
13'b1001001111000,
13'b1001010000011,
13'b1001010000101,
13'b1001010000110,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010000110111,
13'b1010000111000,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001000110,
13'b1010001000111,
13'b1010001001000,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001010110,
13'b1010001010111,
13'b1010001011000,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1010001100101,
13'b1010001100110,
13'b1010001100111,
13'b1010001101000,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010001110111,
13'b1010010000101,
13'b1010010000110,
13'b1011000110101,
13'b1011000110110,
13'b1011000110111,
13'b1011000111000,
13'b1011001000011,
13'b1011001000100,
13'b1011001000101,
13'b1011001000110,
13'b1011001000111,
13'b1011001001000,
13'b1011001010011,
13'b1011001010100,
13'b1011001010101,
13'b1011001010110,
13'b1011001010111,
13'b1011001011000,
13'b1011001100011,
13'b1011001100100,
13'b1011001100101,
13'b1011001100110,
13'b1011001100111,
13'b1011001101000,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011001110111,
13'b1011010000101,
13'b1100000110110,
13'b1100000110111,
13'b1100001000100,
13'b1100001000101,
13'b1100001000110,
13'b1100001000111,
13'b1100001010100,
13'b1100001010101,
13'b1100001010110,
13'b1100001010111,
13'b1100001100101,
13'b1100001100110,
13'b1100001100111,
13'b1100001110101,
13'b1100001110110,
13'b1100001110111: edge_mask_reg_512p3[494] <= 1'b1;
 		default: edge_mask_reg_512p3[494] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[495] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000110,
13'b100000111,
13'b100001000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1100000110,
13'b1100000111,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110110,
13'b100011110111,
13'b101001000111,
13'b101001001000,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110110,
13'b101011110111,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010001000,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000011,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010010,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100000,
13'b1001010100001,
13'b1001010100010,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110000,
13'b1001010110001,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010011,
13'b1010001110011,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000010,
13'b1010010000011,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010000,
13'b1010010010001,
13'b1010010010010,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100000,
13'b1010010100001,
13'b1010010100010,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110000,
13'b1010010110001,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000001,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010010000,
13'b1011010010001,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100000,
13'b1011010100001,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110000,
13'b1011010110001,
13'b1011010110010,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010000,
13'b1100010010001,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010100000,
13'b1100010100001,
13'b1100010100010,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010110000,
13'b1100010110001,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100011000010,
13'b1100011000011,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101010000001,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1101010010000,
13'b1101010010001,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010010101,
13'b1101010100000,
13'b1101010100001,
13'b1101010100010,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010110011,
13'b1101010110100,
13'b1110010000001,
13'b1110010000010,
13'b1110010000011,
13'b1110010000100,
13'b1110010010001,
13'b1110010010010,
13'b1110010010011,
13'b1110010010100,
13'b1110010100001,
13'b1110010100010,
13'b1111010000010,
13'b1111010010010: edge_mask_reg_512p3[496] <= 1'b1;
 		default: edge_mask_reg_512p3[496] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010110,
13'b10010111,
13'b10011000,
13'b10100110,
13'b10100111,
13'b10101000,
13'b10110110,
13'b10110111,
13'b10111000,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11110110,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000110,
13'b100000111,
13'b100001000,
13'b100010110,
13'b100010111,
13'b100011000,
13'b100100110,
13'b100100111,
13'b100101000,
13'b100110110,
13'b100110111,
13'b100111000,
13'b101000110,
13'b101000111,
13'b101001000,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011110110,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1100000110,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100010110,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100110,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b1100110110,
13'b1100110111,
13'b1100111000,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011011001,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011110110,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10100000110,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100010110,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100100111,
13'b10100101000,
13'b10100101001,
13'b10100110111,
13'b10100111000,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011110110,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11100000110,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100100111,
13'b11100101000,
13'b11100101001,
13'b11100111000,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011110110,
13'b100011110111,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100000111,
13'b100100001000,
13'b100100001001,
13'b100100010111,
13'b100100011000,
13'b100100011001,
13'b100100100111,
13'b100100101000,
13'b100100101001,
13'b100100110111,
13'b100100111000,
13'b101001000111,
13'b101001001000,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011110110,
13'b101011110111,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100000111,
13'b101100001000,
13'b101100001001,
13'b101100010111,
13'b101100011000,
13'b101100011001,
13'b101100100111,
13'b101100101000,
13'b101100101001,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011100110,
13'b110011100111,
13'b110011101000,
13'b110011101001,
13'b110011110110,
13'b110011110111,
13'b110011111000,
13'b110011111001,
13'b110100000111,
13'b110100001000,
13'b110100001001,
13'b110100010111,
13'b110100011000,
13'b110100011001,
13'b110100101000,
13'b111001110101,
13'b111001110110,
13'b111001110111,
13'b111010000101,
13'b111010000110,
13'b111010000111,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010011000,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010101000,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111010111000,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011001000,
13'b111011010110,
13'b111011010111,
13'b111011011000,
13'b111011100110,
13'b111011100111,
13'b111011101000,
13'b111011110110,
13'b111011110111,
13'b111011111000,
13'b111100000111,
13'b1000001110100,
13'b1000001110101,
13'b1000001110110,
13'b1000010000100,
13'b1000010000101,
13'b1000010000110,
13'b1000010000111,
13'b1000010010101,
13'b1000010010110,
13'b1000010010111,
13'b1000010100101,
13'b1000010100110,
13'b1000010100111,
13'b1000010110101,
13'b1000010110110,
13'b1000010110111,
13'b1000011000101,
13'b1000011000110,
13'b1000011000111,
13'b1000011010101,
13'b1000011010110,
13'b1000011010111,
13'b1000011011000,
13'b1000011100101,
13'b1000011100110,
13'b1000011100111,
13'b1000011101000,
13'b1000011110110,
13'b1000011110111,
13'b1001001110100,
13'b1001001110101,
13'b1001001110110,
13'b1001010000100,
13'b1001010000101,
13'b1001010000110,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010010111,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010100111,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001010110111,
13'b1001011000101,
13'b1001011000110,
13'b1001011000111,
13'b1001011010101,
13'b1001011010110,
13'b1001011010111,
13'b1001011100101,
13'b1001011100110,
13'b1001011100111,
13'b1001011110101,
13'b1001011110110,
13'b1001011110111,
13'b1001100000110,
13'b1010001110100,
13'b1010001110101,
13'b1010001110110,
13'b1010010000100,
13'b1010010000101,
13'b1010010000110,
13'b1010010010100,
13'b1010010010101,
13'b1010010010110,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010100111,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010010110111,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011000111,
13'b1010011010101,
13'b1010011010110,
13'b1010011010111,
13'b1010011100101,
13'b1010011100110,
13'b1010011100111,
13'b1010011110101,
13'b1010011110110,
13'b1010011110111,
13'b1010100000101,
13'b1010100000110,
13'b1011001110011,
13'b1011001110100,
13'b1011001110101,
13'b1011001110110,
13'b1011010000010,
13'b1011010000011,
13'b1011010000100,
13'b1011010000101,
13'b1011010000110,
13'b1011010010010,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010010110,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010100110,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011010110110,
13'b1011011000100,
13'b1011011000101,
13'b1011011000110,
13'b1011011000111,
13'b1011011010100,
13'b1011011010101,
13'b1011011010110,
13'b1011011010111,
13'b1011011100100,
13'b1011011100101,
13'b1011011100110,
13'b1011011100111,
13'b1011011110100,
13'b1011011110101,
13'b1011011110110,
13'b1011011110111,
13'b1011100000101,
13'b1011100000110,
13'b1100001110011,
13'b1100001110100,
13'b1100001110101,
13'b1100010000001,
13'b1100010000010,
13'b1100010000011,
13'b1100010000100,
13'b1100010000101,
13'b1100010010001,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010010110,
13'b1100010100001,
13'b1100010100010,
13'b1100010100011,
13'b1100010100100,
13'b1100010100101,
13'b1100010100110,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100010110101,
13'b1100010110110,
13'b1100011000010,
13'b1100011000011,
13'b1100011000100,
13'b1100011000101,
13'b1100011000110,
13'b1100011010011,
13'b1100011010100,
13'b1100011010101,
13'b1100011010110,
13'b1100011100011,
13'b1100011100100,
13'b1100011100101,
13'b1100011100110,
13'b1100011110100,
13'b1100011110101,
13'b1100011110110,
13'b1100100000101,
13'b1101001110011,
13'b1101001110100,
13'b1101001110101,
13'b1101010000001,
13'b1101010000010,
13'b1101010000011,
13'b1101010000100,
13'b1101010000101,
13'b1101010010001,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010010101,
13'b1101010100001,
13'b1101010100010,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010110010,
13'b1101010110011,
13'b1101010110100,
13'b1101010110101,
13'b1101010110110,
13'b1101011000010,
13'b1101011000011,
13'b1101011000100,
13'b1101011000101,
13'b1101011000110,
13'b1101011010010,
13'b1101011010011,
13'b1101011010100,
13'b1101011010101,
13'b1101011010110,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011100101,
13'b1101011100110,
13'b1101011110011,
13'b1101011110100,
13'b1101011110101,
13'b1101011110110,
13'b1101100000101,
13'b1110010000001,
13'b1110010000010,
13'b1110010000011,
13'b1110010000100,
13'b1110010010010,
13'b1110010010011,
13'b1110010010100,
13'b1110010010101,
13'b1110010100010,
13'b1110010100011,
13'b1110010100100,
13'b1110010100101,
13'b1110010110010,
13'b1110010110011,
13'b1110010110100,
13'b1110010110101,
13'b1110011000010,
13'b1110011000011,
13'b1110011000100,
13'b1110011000101,
13'b1110011000110,
13'b1110011010010,
13'b1110011010011,
13'b1110011010100,
13'b1110011010101,
13'b1110011010110,
13'b1110011100010,
13'b1110011100011,
13'b1110011100100,
13'b1110011100101,
13'b1110011100110,
13'b1110011110011,
13'b1110011110100,
13'b1110011110101,
13'b1110011110110,
13'b1111010000010,
13'b1111010010010,
13'b1111010010011,
13'b1111010100010,
13'b1111010100011,
13'b1111010100100,
13'b1111010110010,
13'b1111010110011,
13'b1111010110100,
13'b1111011000010,
13'b1111011000011,
13'b1111011000100,
13'b1111011010010,
13'b1111011010011,
13'b1111011010100,
13'b1111011010101,
13'b1111011100011,
13'b1111011100100,
13'b1111011100101,
13'b1111011110011,
13'b1111011110100: edge_mask_reg_512p3[497] <= 1'b1;
 		default: edge_mask_reg_512p3[497] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10001010101,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010101,
13'b100001010110,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000101,
13'b101001000110,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000101,
13'b110001000110,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100011,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100011,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000100010,
13'b1001000100011,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100010,
13'b1010000100011,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000100001,
13'b1101000000000,
13'b1101000000001,
13'b1101000000010,
13'b1101000000011,
13'b1101000010000,
13'b1101000010001,
13'b1101000010010,
13'b1101000010011,
13'b1110000000000,
13'b1110000000001,
13'b1110000010000: edge_mask_reg_512p3[498] <= 1'b1;
 		default: edge_mask_reg_512p3[498] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[499] <= 1'b0;
 	endcase

    case({x,y,z})
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b11001000100,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001110101,
13'b11001110110,
13'b100000110100,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100001000100,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b101000100011,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001110101,
13'b101001110110,
13'b110000100010,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001100101,
13'b110001100110,
13'b111000010001,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b1000000010000,
13'b1000000010001,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100001,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000011,
13'b1000001000100,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000100000,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1101000000000,
13'b1101000010000,
13'b1101000010001,
13'b1101000100000,
13'b1101000100001,
13'b1101000100010,
13'b1101000110000,
13'b1101000110001,
13'b1101000110010,
13'b1101001000000,
13'b1110000010000,
13'b1110000100000,
13'b1110000110000: edge_mask_reg_512p3[500] <= 1'b1;
 		default: edge_mask_reg_512p3[500] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[501] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[502] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[503] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100101,
13'b10100110,
13'b10100111,
13'b10110101,
13'b10110110,
13'b10110111,
13'b11000101,
13'b11000110,
13'b11000111,
13'b11001000,
13'b11010101,
13'b11010110,
13'b11010111,
13'b11011000,
13'b11100101,
13'b11100110,
13'b11100111,
13'b11101000,
13'b11110101,
13'b11110110,
13'b11110111,
13'b11111000,
13'b100000101,
13'b100000110,
13'b100000111,
13'b100010101,
13'b100010110,
13'b100010111,
13'b100100101,
13'b100100110,
13'b100100111,
13'b100110101,
13'b100110110,
13'b100110111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1001111000,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010001000,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b1010011000,
13'b1010100101,
13'b1010100110,
13'b1010100111,
13'b1010101000,
13'b1010110101,
13'b1010110110,
13'b1010110111,
13'b1010111000,
13'b1011000101,
13'b1011000110,
13'b1011000111,
13'b1011001000,
13'b1011010101,
13'b1011010110,
13'b1011010111,
13'b1011011000,
13'b1011100101,
13'b1011100110,
13'b1011100111,
13'b1011101000,
13'b1011110101,
13'b1011110110,
13'b1011110111,
13'b1100000101,
13'b1100000110,
13'b1100000111,
13'b1100010101,
13'b1100010110,
13'b1100010111,
13'b1100100101,
13'b1100100110,
13'b1100100111,
13'b10001010110,
13'b10001010111,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10001111000,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010001000,
13'b10010010100,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b10010011000,
13'b10010100100,
13'b10010100101,
13'b10010100110,
13'b10010100111,
13'b10010101000,
13'b10010110100,
13'b10010110101,
13'b10010110110,
13'b10010110111,
13'b10010111000,
13'b10011000100,
13'b10011000101,
13'b10011000110,
13'b10011000111,
13'b10011001000,
13'b10011010100,
13'b10011010101,
13'b10011010110,
13'b10011010111,
13'b10011011000,
13'b10011100100,
13'b10011100101,
13'b10011100110,
13'b10011100111,
13'b10011101000,
13'b10011110100,
13'b10011110101,
13'b10011110110,
13'b10011110111,
13'b10100000100,
13'b10100000101,
13'b10100000110,
13'b10100000111,
13'b10100010100,
13'b10100010101,
13'b10100010110,
13'b10100010111,
13'b10100100101,
13'b10100100110,
13'b10100100111,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010110100,
13'b11010110101,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11011000100,
13'b11011000101,
13'b11011000110,
13'b11011000111,
13'b11011001000,
13'b11011010100,
13'b11011010101,
13'b11011010110,
13'b11011010111,
13'b11011011000,
13'b11011100100,
13'b11011100101,
13'b11011100110,
13'b11011100111,
13'b11011101000,
13'b11011110100,
13'b11011110101,
13'b11011110110,
13'b11011110111,
13'b11100000100,
13'b11100000101,
13'b11100000110,
13'b11100000111,
13'b11100010100,
13'b11100010101,
13'b11100010110,
13'b11100010111,
13'b11100100101,
13'b11100100110,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010110100,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100011000100,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011010100,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011100100,
13'b100011100101,
13'b100011100110,
13'b100011100111,
13'b100011101000,
13'b100011110100,
13'b100011110101,
13'b100011110110,
13'b100011110111,
13'b100100000100,
13'b100100000101,
13'b100100000110,
13'b100100000111,
13'b100100010100,
13'b100100010101,
13'b100100010110,
13'b100100010111,
13'b100100100101,
13'b100100100110,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011100100,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011110100,
13'b101011110101,
13'b101011110110,
13'b101011110111,
13'b101100000100,
13'b101100000101,
13'b101100000110,
13'b101100000111,
13'b101100010100,
13'b101100010101,
13'b101100010110,
13'b101100100101,
13'b101100100110,
13'b110001100110,
13'b110001100111,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011100011,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b110011110100,
13'b110011110101,
13'b110011110110,
13'b110011110111,
13'b110100000100,
13'b110100000101,
13'b110100000110,
13'b110100010101,
13'b110100010110,
13'b111010000101,
13'b111010000110,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b111011110100,
13'b111011110101,
13'b1000010010100,
13'b1000010010101,
13'b1000010010110,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011110011,
13'b1000011110100,
13'b1001010010011,
13'b1001010010100,
13'b1001010010101,
13'b1001010010110,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010100110,
13'b1001010110010,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001010110110,
13'b1001011000010,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011000110,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101,
13'b1001011110011,
13'b1001011110100,
13'b1010010000100,
13'b1010010000101,
13'b1010010010011,
13'b1010010010100,
13'b1010010010101,
13'b1010010100011,
13'b1010010100100,
13'b1010010100101,
13'b1010010100110,
13'b1010010110010,
13'b1010010110011,
13'b1010010110100,
13'b1010010110101,
13'b1010010110110,
13'b1010011000010,
13'b1010011000011,
13'b1010011000100,
13'b1010011000101,
13'b1010011000110,
13'b1010011010010,
13'b1010011010011,
13'b1010011010100,
13'b1010011010101,
13'b1010011100010,
13'b1010011100011,
13'b1010011100100,
13'b1010011100101,
13'b1010011110010,
13'b1010011110011,
13'b1010011110100,
13'b1011010000100,
13'b1011010010011,
13'b1011010010100,
13'b1011010010101,
13'b1011010100010,
13'b1011010100011,
13'b1011010100100,
13'b1011010100101,
13'b1011010110010,
13'b1011010110011,
13'b1011010110100,
13'b1011010110101,
13'b1011011000001,
13'b1011011000010,
13'b1011011000011,
13'b1011011000100,
13'b1011011000101,
13'b1011011010001,
13'b1011011010010,
13'b1011011010011,
13'b1011011010100,
13'b1011011010101,
13'b1011011100010,
13'b1011011100011,
13'b1011011100100,
13'b1011011110010,
13'b1011011110011,
13'b1011011110100,
13'b1100010000100,
13'b1100010010010,
13'b1100010010011,
13'b1100010010100,
13'b1100010010101,
13'b1100010100001,
13'b1100010100010,
13'b1100010100011,
13'b1100010100100,
13'b1100010110000,
13'b1100010110001,
13'b1100010110010,
13'b1100010110011,
13'b1100010110100,
13'b1100010110101,
13'b1100011000000,
13'b1100011000001,
13'b1100011000010,
13'b1100011000011,
13'b1100011000100,
13'b1100011000101,
13'b1100011010000,
13'b1100011010001,
13'b1100011010010,
13'b1100011010011,
13'b1100011010100,
13'b1100011100000,
13'b1100011100001,
13'b1100011100010,
13'b1100011100011,
13'b1100011100100,
13'b1100011110010,
13'b1100011110011,
13'b1101010010010,
13'b1101010010011,
13'b1101010010100,
13'b1101010100001,
13'b1101010100010,
13'b1101010100011,
13'b1101010100100,
13'b1101010100101,
13'b1101010110000,
13'b1101010110001,
13'b1101010110010,
13'b1101010110011,
13'b1101010110100,
13'b1101010110101,
13'b1101011000000,
13'b1101011000001,
13'b1101011000010,
13'b1101011000011,
13'b1101011000100,
13'b1101011010000,
13'b1101011010001,
13'b1101011010010,
13'b1101011010011,
13'b1101011010100,
13'b1101011100000,
13'b1101011100001,
13'b1101011100010,
13'b1101011100011,
13'b1101011100100,
13'b1101011110000,
13'b1101011110001,
13'b1101011110010,
13'b1101011110011,
13'b1110010010011,
13'b1110010010100,
13'b1110010100001,
13'b1110010100010,
13'b1110010100011,
13'b1110010100100,
13'b1110010110000,
13'b1110010110001,
13'b1110010110010,
13'b1110010110011,
13'b1110010110100,
13'b1110011000000,
13'b1110011000001,
13'b1110011000010,
13'b1110011000011,
13'b1110011000100,
13'b1110011010000,
13'b1110011010001,
13'b1110011010010,
13'b1110011010011,
13'b1110011010100,
13'b1110011100000,
13'b1110011100001,
13'b1110011100010,
13'b1110011100011,
13'b1110011100100,
13'b1110011110000,
13'b1110011110001,
13'b1110011110010,
13'b1110011110011,
13'b1111010100001,
13'b1111010100010,
13'b1111010110001,
13'b1111010110010,
13'b1111011000000,
13'b1111011000001,
13'b1111011000010,
13'b1111011010000,
13'b1111011010001,
13'b1111011010010,
13'b1111011100000,
13'b1111011100001,
13'b1111011110000: edge_mask_reg_512p3[504] <= 1'b1;
 		default: edge_mask_reg_512p3[504] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b100111000,
13'b100111001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100100111,
13'b1100101000,
13'b1100101001,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100010111,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b10100101001,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011110111,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100000111,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100010111,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b11100101000,
13'b11100101001,
13'b100001111000,
13'b100001111001,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b100100101000,
13'b100100101001,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b101100011000,
13'b101100011001,
13'b110010011000,
13'b110010011001,
13'b110010101000,
13'b110010101001,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011101000,
13'b110011101001,
13'b110011101010,
13'b110011111000,
13'b110011111001,
13'b110100001000,
13'b110100001001,
13'b111010101000,
13'b111010101001,
13'b111010111000,
13'b111010111001,
13'b111010111010,
13'b111011001000,
13'b111011001001,
13'b111011001010,
13'b111011010111,
13'b111011011000,
13'b111011011001,
13'b111011011010,
13'b111011101000,
13'b111011101001,
13'b1000010101000,
13'b1000010101001,
13'b1000010111000,
13'b1000010111001,
13'b1000010111010,
13'b1000011000111,
13'b1000011001000,
13'b1000011001001,
13'b1000011001010,
13'b1000011010111,
13'b1000011011000,
13'b1000011011001,
13'b1000011100111,
13'b1000011101000,
13'b1000011101001,
13'b1001010101000,
13'b1001010101001,
13'b1001010111000,
13'b1001010111001,
13'b1001010111010,
13'b1001011000111,
13'b1001011001000,
13'b1001011001001,
13'b1001011001010,
13'b1001011010111,
13'b1001011011000,
13'b1001011011001,
13'b1001011100111,
13'b1001011101000,
13'b1001011101001,
13'b1010010101000,
13'b1010010101001,
13'b1010010111000,
13'b1010010111001,
13'b1010010111010,
13'b1010011000111,
13'b1010011001000,
13'b1010011001001,
13'b1010011001010,
13'b1010011010111,
13'b1010011011000,
13'b1010011011001,
13'b1010011100111,
13'b1010011101000,
13'b1010011101001,
13'b1011010101000,
13'b1011010101001,
13'b1011010111000,
13'b1011010111001,
13'b1011010111010,
13'b1011011000111,
13'b1011011001000,
13'b1011011001001,
13'b1011011001010,
13'b1011011010111,
13'b1011011011000,
13'b1011011011001,
13'b1011011100111,
13'b1011011101000,
13'b1011011101001,
13'b1100010101000,
13'b1100010101001,
13'b1100010110111,
13'b1100010111000,
13'b1100010111001,
13'b1100010111010,
13'b1100011000111,
13'b1100011001000,
13'b1100011001001,
13'b1100011001010,
13'b1100011010111,
13'b1100011011000,
13'b1100011011001,
13'b1100011100111,
13'b1100011101000,
13'b1100011101001,
13'b1101010101000,
13'b1101010101001,
13'b1101010110111,
13'b1101010111000,
13'b1101010111001,
13'b1101010111010,
13'b1101011000111,
13'b1101011001000,
13'b1101011001001,
13'b1101011001010,
13'b1101011010110,
13'b1101011010111,
13'b1101011011000,
13'b1101011011001,
13'b1101011011010,
13'b1101011100110,
13'b1101011100111,
13'b1101011101000,
13'b1101011101001,
13'b1110010101001,
13'b1110010110111,
13'b1110010111000,
13'b1110010111001,
13'b1110010111010,
13'b1110011000111,
13'b1110011001000,
13'b1110011001001,
13'b1110011001010,
13'b1110011010111,
13'b1110011011000,
13'b1110011011001,
13'b1110011011010,
13'b1110011100111,
13'b1110011101000,
13'b1110011101001,
13'b1111010110111,
13'b1111010111000,
13'b1111010111001,
13'b1111011000110,
13'b1111011000111,
13'b1111011001000,
13'b1111011001001,
13'b1111011010110,
13'b1111011010111,
13'b1111011011000,
13'b1111011011001: edge_mask_reg_512p3[505] <= 1'b1;
 		default: edge_mask_reg_512p3[505] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10110111,
13'b10111000,
13'b10111001,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11100111,
13'b11101000,
13'b11101001,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010110111,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10011000111,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011011000,
13'b10011011001,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000100,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010011,
13'b11010010100,
13'b11010010101,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100100,
13'b11010100101,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011011000,
13'b11011011001,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011011000,
13'b100011011001,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000101011,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101000111011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001001011,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001011011,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010010001,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010110100,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011001000,
13'b101011001001,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110000111010,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111001,
13'b110001111010,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001001,
13'b110010001010,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010011001,
13'b110010011010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010101001,
13'b110010110011,
13'b110010110100,
13'b110010111001,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000101000,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111000111000,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001001000,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001100111,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010100011,
13'b111010100100,
13'b1000000010100,
13'b1000000010101,
13'b1000000010110,
13'b1000000010111,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000100110,
13'b1000000100111,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000000110110,
13'b1000000110111,
13'b1000001000001,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001000110,
13'b1000001000111,
13'b1000001010001,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001010110,
13'b1000001010111,
13'b1000001100001,
13'b1000001100010,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001100110,
13'b1000001110001,
13'b1000001110010,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000010000001,
13'b1000010000010,
13'b1000010000011,
13'b1000010000100,
13'b1001000010100,
13'b1001000010101,
13'b1001000010110,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000100110,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001000110110,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001000110,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001010110,
13'b1001001100001,
13'b1001001100010,
13'b1001001100011,
13'b1001001100100,
13'b1001001100101,
13'b1001001110001,
13'b1001001110010,
13'b1001001110011,
13'b1010000010100,
13'b1010000010101,
13'b1010000010110,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000100101,
13'b1010000100110,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010000110101,
13'b1010000110110,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001000101,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001100010,
13'b1010001100011,
13'b1011000100011,
13'b1011000100100,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001010010,
13'b1011001010011: edge_mask_reg_512p3[506] <= 1'b1;
 		default: edge_mask_reg_512p3[506] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010101,
13'b10010110,
13'b10010111,
13'b10100110,
13'b10100111,
13'b1001100101,
13'b1001100110,
13'b1001100111,
13'b1001101000,
13'b1001110101,
13'b1001110110,
13'b1001110111,
13'b1010000101,
13'b1010000110,
13'b1010000111,
13'b1010010101,
13'b1010010110,
13'b1010010111,
13'b10001010101,
13'b10001010110,
13'b10001010111,
13'b10001011000,
13'b10001100101,
13'b10001100110,
13'b10001100111,
13'b10001101000,
13'b10001110101,
13'b10001110110,
13'b10001110111,
13'b10010000101,
13'b10010000110,
13'b10010000111,
13'b10010010101,
13'b10010010110,
13'b10010010111,
13'b11001000101,
13'b11001000110,
13'b11001000111,
13'b11001001000,
13'b11001010101,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001100101,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001110101,
13'b11001110110,
13'b11001110111,
13'b11010000101,
13'b11010000110,
13'b11010000111,
13'b11010010110,
13'b11010010111,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010010110,
13'b100010010111,
13'b101000100100,
13'b101000100101,
13'b101000100110,
13'b101000100111,
13'b101000101000,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010010110,
13'b101010010111,
13'b110000100011,
13'b110000100100,
13'b110000100101,
13'b110000100110,
13'b110000100111,
13'b110000101000,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110010000110,
13'b110010000111,
13'b111000010010,
13'b111000010011,
13'b111000010100,
13'b111000010101,
13'b111000010110,
13'b111000010111,
13'b111000100010,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000100110,
13'b111000100111,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111000110111,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001010111,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b1000000010010,
13'b1000000010011,
13'b1000000010100,
13'b1000000010101,
13'b1000000100010,
13'b1000000100011,
13'b1000000100100,
13'b1000000100101,
13'b1000000110010,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001100011,
13'b1000001100100,
13'b1001000010000,
13'b1001000010001,
13'b1001000010010,
13'b1001000010011,
13'b1001000010100,
13'b1001000100001,
13'b1001000100010,
13'b1001000100011,
13'b1001000100100,
13'b1001000100101,
13'b1001000110001,
13'b1001000110010,
13'b1001000110011,
13'b1001000110100,
13'b1001000110101,
13'b1001001000001,
13'b1001001000010,
13'b1001001000011,
13'b1001001000100,
13'b1001001000101,
13'b1001001010001,
13'b1001001010010,
13'b1001001010011,
13'b1001001010100,
13'b1001001010101,
13'b1001001100011,
13'b1001001100100,
13'b1010000000000,
13'b1010000000001,
13'b1010000000010,
13'b1010000000011,
13'b1010000000100,
13'b1010000010000,
13'b1010000010001,
13'b1010000010010,
13'b1010000010011,
13'b1010000010100,
13'b1010000100000,
13'b1010000100001,
13'b1010000100010,
13'b1010000100011,
13'b1010000100100,
13'b1010000110000,
13'b1010000110001,
13'b1010000110010,
13'b1010000110011,
13'b1010000110100,
13'b1010001000000,
13'b1010001000001,
13'b1010001000010,
13'b1010001000011,
13'b1010001000100,
13'b1010001010000,
13'b1010001010001,
13'b1010001010010,
13'b1010001010011,
13'b1010001010100,
13'b1010001010101,
13'b1010001100000,
13'b1010001100001,
13'b1010001100010,
13'b1010001100011,
13'b1010001100100,
13'b1011000000000,
13'b1011000000001,
13'b1011000000010,
13'b1011000000011,
13'b1011000010000,
13'b1011000010001,
13'b1011000010010,
13'b1011000010011,
13'b1011000100000,
13'b1011000100001,
13'b1011000100010,
13'b1011000100011,
13'b1011000110000,
13'b1011000110001,
13'b1011000110010,
13'b1011000110011,
13'b1011000110100,
13'b1011001000000,
13'b1011001000001,
13'b1011001000010,
13'b1011001000011,
13'b1011001000100,
13'b1011001010000,
13'b1011001010001,
13'b1011001010010,
13'b1011001010011,
13'b1011001010100,
13'b1011001100000,
13'b1011001100001,
13'b1011001100010,
13'b1011001100011,
13'b1011001100100,
13'b1100000000000,
13'b1100000000001,
13'b1100000000010,
13'b1100000000011,
13'b1100000010000,
13'b1100000010001,
13'b1100000010010,
13'b1100000010011,
13'b1100000100000,
13'b1100000100001,
13'b1100000100010,
13'b1100000100011,
13'b1100000110000,
13'b1100000110001,
13'b1100000110010,
13'b1100000110011,
13'b1100001000000,
13'b1100001000001,
13'b1100001000010,
13'b1100001000011,
13'b1100001010000,
13'b1100001010001,
13'b1100001010010,
13'b1100001010011,
13'b1100001100000,
13'b1100001100001,
13'b1100001100010,
13'b1101001000000,
13'b1101001000010,
13'b1101001000011,
13'b1101001010000,
13'b1101001010010,
13'b1101001010011,
13'b1101001100000: edge_mask_reg_512p3[507] <= 1'b1;
 		default: edge_mask_reg_512p3[507] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[508] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b11110111,
13'b11111000,
13'b11111001,
13'b11111010,
13'b100000111,
13'b100001000,
13'b100001001,
13'b100010111,
13'b100011000,
13'b100011001,
13'b100100111,
13'b100101000,
13'b100101001,
13'b1001100111,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011010111,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b1011011011,
13'b1011100111,
13'b1011101000,
13'b1011101001,
13'b1011101010,
13'b1011110111,
13'b1011111000,
13'b1011111001,
13'b1011111010,
13'b1100000111,
13'b1100001000,
13'b1100001001,
13'b1100001010,
13'b1100010111,
13'b1100011000,
13'b1100011001,
13'b1100011010,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010101100,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b10011011011,
13'b10011100111,
13'b10011101000,
13'b10011101001,
13'b10011101010,
13'b10011101011,
13'b10011110111,
13'b10011111000,
13'b10011111001,
13'b10011111010,
13'b10100000111,
13'b10100001000,
13'b10100001001,
13'b10100001010,
13'b10100011000,
13'b10100011001,
13'b10100011010,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100010,
13'b11001100011,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110010,
13'b11001110011,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000010,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010010,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010110110,
13'b11010110111,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011000111,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011010111,
13'b11011011000,
13'b11011011001,
13'b11011011010,
13'b11011011011,
13'b11011100111,
13'b11011101000,
13'b11011101001,
13'b11011101010,
13'b11011101011,
13'b11011111000,
13'b11011111001,
13'b11011111010,
13'b11100001000,
13'b11100001001,
13'b11100001010,
13'b11100011000,
13'b11100011001,
13'b11100011010,
13'b100000111001,
13'b100000111010,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010101,
13'b100001010110,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100010,
13'b100010100011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010110010,
13'b100010110101,
13'b100010110110,
13'b100010110111,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011000101,
13'b100011000110,
13'b100011000111,
13'b100011001000,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011010101,
13'b100011010110,
13'b100011010111,
13'b100011011000,
13'b100011011001,
13'b100011011010,
13'b100011011011,
13'b100011100111,
13'b100011101000,
13'b100011101001,
13'b100011101010,
13'b100011111000,
13'b100011111001,
13'b100011111010,
13'b100100001000,
13'b100100001001,
13'b100100001010,
13'b100100011000,
13'b100100011001,
13'b100100011010,
13'b101001001001,
13'b101001001010,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001011001,
13'b101001011010,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100010,
13'b101010100011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010101011,
13'b101010110010,
13'b101010110011,
13'b101010110100,
13'b101010110101,
13'b101010110110,
13'b101010110111,
13'b101010111000,
13'b101010111001,
13'b101010111010,
13'b101011000010,
13'b101011000011,
13'b101011000100,
13'b101011000101,
13'b101011000110,
13'b101011000111,
13'b101011001000,
13'b101011001001,
13'b101011001010,
13'b101011010100,
13'b101011010101,
13'b101011010110,
13'b101011010111,
13'b101011011000,
13'b101011011001,
13'b101011011010,
13'b101011100101,
13'b101011100110,
13'b101011100111,
13'b101011101000,
13'b101011101001,
13'b101011101010,
13'b101011111000,
13'b101011111001,
13'b101011111010,
13'b101100001000,
13'b101100001001,
13'b101100001010,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111010,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001001,
13'b110010001010,
13'b110010010001,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011000,
13'b110010011001,
13'b110010011010,
13'b110010100001,
13'b110010100010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b110010101000,
13'b110010101001,
13'b110010101010,
13'b110010110001,
13'b110010110010,
13'b110010110011,
13'b110010110100,
13'b110010110101,
13'b110010110110,
13'b110010110111,
13'b110010111000,
13'b110010111001,
13'b110010111010,
13'b110011000001,
13'b110011000010,
13'b110011000011,
13'b110011000100,
13'b110011000101,
13'b110011000110,
13'b110011000111,
13'b110011001000,
13'b110011001001,
13'b110011001010,
13'b110011010001,
13'b110011010010,
13'b110011010011,
13'b110011010100,
13'b110011010101,
13'b110011010110,
13'b110011010111,
13'b110011011000,
13'b110011011001,
13'b110011011010,
13'b110011100100,
13'b110011100101,
13'b110011100110,
13'b110011100111,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111010000001,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010010001,
13'b111010010010,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010010111,
13'b111010100001,
13'b111010100010,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b111010100110,
13'b111010100111,
13'b111010110001,
13'b111010110010,
13'b111010110011,
13'b111010110100,
13'b111010110101,
13'b111010110110,
13'b111010110111,
13'b111011000001,
13'b111011000010,
13'b111011000011,
13'b111011000100,
13'b111011000101,
13'b111011000110,
13'b111011000111,
13'b111011010001,
13'b111011010010,
13'b111011010011,
13'b111011010100,
13'b111011010101,
13'b111011010110,
13'b111011010111,
13'b111011100011,
13'b111011100100,
13'b111011100101,
13'b111011100110,
13'b1000001100100,
13'b1000001110100,
13'b1000001110101,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010010,
13'b1000010010011,
13'b1000010010100,
13'b1000010010101,
13'b1000010100001,
13'b1000010100010,
13'b1000010100011,
13'b1000010100100,
13'b1000010100101,
13'b1000010100110,
13'b1000010110001,
13'b1000010110010,
13'b1000010110011,
13'b1000010110100,
13'b1000010110101,
13'b1000010110110,
13'b1000011000001,
13'b1000011000010,
13'b1000011000011,
13'b1000011000100,
13'b1000011000101,
13'b1000011000110,
13'b1000011010001,
13'b1000011010010,
13'b1000011010011,
13'b1000011010100,
13'b1000011010101,
13'b1000011010110,
13'b1000011100011,
13'b1000011100100,
13'b1000011100101,
13'b1000011100110,
13'b1001010010100,
13'b1001010100011,
13'b1001010100100,
13'b1001010100101,
13'b1001010110011,
13'b1001010110100,
13'b1001010110101,
13'b1001011000011,
13'b1001011000100,
13'b1001011000101,
13'b1001011010010,
13'b1001011010011,
13'b1001011010100,
13'b1001011010101,
13'b1001011100011,
13'b1001011100100,
13'b1001011100101: edge_mask_reg_512p3[509] <= 1'b1;
 		default: edge_mask_reg_512p3[509] <= 1'b0;
 	endcase

    case({x,y,z})
13'b10010111,
13'b10011000,
13'b10011001,
13'b10011010,
13'b10011011,
13'b10100111,
13'b10101000,
13'b10101001,
13'b10101010,
13'b10101011,
13'b10110111,
13'b10111000,
13'b10111001,
13'b10111010,
13'b11000111,
13'b11001000,
13'b11001001,
13'b11001010,
13'b11010111,
13'b11011000,
13'b11011001,
13'b11011010,
13'b11100111,
13'b11101000,
13'b11101001,
13'b11101010,
13'b1001101000,
13'b1001101001,
13'b1001101010,
13'b1001101011,
13'b1001101100,
13'b1001110111,
13'b1001111000,
13'b1001111001,
13'b1001111010,
13'b1001111011,
13'b1001111100,
13'b1010000111,
13'b1010001000,
13'b1010001001,
13'b1010001010,
13'b1010001011,
13'b1010001100,
13'b1010010111,
13'b1010011000,
13'b1010011001,
13'b1010011010,
13'b1010011011,
13'b1010011100,
13'b1010100111,
13'b1010101000,
13'b1010101001,
13'b1010101010,
13'b1010101011,
13'b1010110111,
13'b1010111000,
13'b1010111001,
13'b1010111010,
13'b1010111011,
13'b1011000111,
13'b1011001000,
13'b1011001001,
13'b1011001010,
13'b1011001011,
13'b1011011000,
13'b1011011001,
13'b1011011010,
13'b10001010111,
13'b10001011000,
13'b10001011001,
13'b10001011010,
13'b10001011011,
13'b10001100111,
13'b10001101000,
13'b10001101001,
13'b10001101010,
13'b10001101011,
13'b10001101100,
13'b10001110111,
13'b10001111000,
13'b10001111001,
13'b10001111010,
13'b10001111011,
13'b10001111100,
13'b10010000111,
13'b10010001000,
13'b10010001001,
13'b10010001010,
13'b10010001011,
13'b10010001100,
13'b10010010111,
13'b10010011000,
13'b10010011001,
13'b10010011010,
13'b10010011011,
13'b10010011100,
13'b10010100111,
13'b10010101000,
13'b10010101001,
13'b10010101010,
13'b10010101011,
13'b10010111000,
13'b10010111001,
13'b10010111010,
13'b10010111011,
13'b10011001000,
13'b10011001001,
13'b10011001010,
13'b10011001011,
13'b10011011000,
13'b10011011001,
13'b10011011010,
13'b11001000111,
13'b11001001000,
13'b11001001001,
13'b11001001010,
13'b11001001011,
13'b11001010110,
13'b11001010111,
13'b11001011000,
13'b11001011001,
13'b11001011010,
13'b11001011011,
13'b11001100010,
13'b11001100011,
13'b11001100110,
13'b11001100111,
13'b11001101000,
13'b11001101001,
13'b11001101010,
13'b11001101011,
13'b11001110010,
13'b11001110011,
13'b11001110110,
13'b11001110111,
13'b11001111000,
13'b11001111001,
13'b11001111010,
13'b11001111011,
13'b11010000010,
13'b11010000110,
13'b11010000111,
13'b11010001000,
13'b11010001001,
13'b11010001010,
13'b11010001011,
13'b11010010010,
13'b11010010110,
13'b11010010111,
13'b11010011000,
13'b11010011001,
13'b11010011010,
13'b11010011011,
13'b11010100110,
13'b11010100111,
13'b11010101000,
13'b11010101001,
13'b11010101010,
13'b11010101011,
13'b11010111000,
13'b11010111001,
13'b11010111010,
13'b11010111011,
13'b11011001000,
13'b11011001001,
13'b11011001010,
13'b11011001011,
13'b11011011001,
13'b11011011010,
13'b100000110101,
13'b100000110110,
13'b100000110111,
13'b100000111000,
13'b100000111001,
13'b100000111010,
13'b100000111011,
13'b100001000001,
13'b100001000010,
13'b100001000101,
13'b100001000110,
13'b100001000111,
13'b100001001000,
13'b100001001001,
13'b100001001010,
13'b100001001011,
13'b100001010001,
13'b100001010010,
13'b100001010011,
13'b100001010101,
13'b100001010110,
13'b100001010111,
13'b100001011000,
13'b100001011001,
13'b100001011010,
13'b100001011011,
13'b100001100001,
13'b100001100010,
13'b100001100011,
13'b100001100100,
13'b100001100101,
13'b100001100110,
13'b100001100111,
13'b100001101000,
13'b100001101001,
13'b100001101010,
13'b100001101011,
13'b100001110001,
13'b100001110010,
13'b100001110011,
13'b100001110100,
13'b100001110101,
13'b100001110110,
13'b100001110111,
13'b100001111000,
13'b100001111001,
13'b100001111010,
13'b100001111011,
13'b100010000010,
13'b100010000011,
13'b100010000100,
13'b100010000101,
13'b100010000110,
13'b100010000111,
13'b100010001000,
13'b100010001001,
13'b100010001010,
13'b100010001011,
13'b100010010010,
13'b100010010011,
13'b100010010100,
13'b100010010101,
13'b100010010110,
13'b100010010111,
13'b100010011000,
13'b100010011001,
13'b100010011010,
13'b100010011011,
13'b100010100100,
13'b100010100101,
13'b100010100110,
13'b100010100111,
13'b100010101000,
13'b100010101001,
13'b100010101010,
13'b100010101011,
13'b100010111000,
13'b100010111001,
13'b100010111010,
13'b100010111011,
13'b100011001001,
13'b100011001010,
13'b100011001011,
13'b100011011001,
13'b100011011010,
13'b101000100101,
13'b101000101000,
13'b101000101001,
13'b101000101010,
13'b101000110001,
13'b101000110010,
13'b101000110011,
13'b101000110100,
13'b101000110101,
13'b101000110110,
13'b101000110111,
13'b101000111000,
13'b101000111001,
13'b101000111010,
13'b101001000001,
13'b101001000010,
13'b101001000011,
13'b101001000100,
13'b101001000101,
13'b101001000110,
13'b101001000111,
13'b101001001000,
13'b101001001001,
13'b101001001010,
13'b101001010001,
13'b101001010010,
13'b101001010011,
13'b101001010100,
13'b101001010101,
13'b101001010110,
13'b101001010111,
13'b101001011000,
13'b101001011001,
13'b101001011010,
13'b101001100001,
13'b101001100010,
13'b101001100011,
13'b101001100100,
13'b101001100101,
13'b101001100110,
13'b101001100111,
13'b101001101000,
13'b101001101001,
13'b101001101010,
13'b101001101011,
13'b101001110001,
13'b101001110010,
13'b101001110011,
13'b101001110100,
13'b101001110101,
13'b101001110110,
13'b101001110111,
13'b101001111000,
13'b101001111001,
13'b101001111010,
13'b101001111011,
13'b101010000001,
13'b101010000010,
13'b101010000011,
13'b101010000100,
13'b101010000101,
13'b101010000110,
13'b101010000111,
13'b101010001000,
13'b101010001001,
13'b101010001010,
13'b101010001011,
13'b101010010010,
13'b101010010011,
13'b101010010100,
13'b101010010101,
13'b101010010110,
13'b101010010111,
13'b101010011000,
13'b101010011001,
13'b101010011010,
13'b101010011011,
13'b101010100100,
13'b101010100101,
13'b101010100110,
13'b101010100111,
13'b101010101000,
13'b101010101001,
13'b101010101010,
13'b101010111001,
13'b101010111010,
13'b110000100100,
13'b110000100101,
13'b110000101000,
13'b110000101001,
13'b110000110001,
13'b110000110010,
13'b110000110011,
13'b110000110100,
13'b110000110101,
13'b110000110110,
13'b110000110111,
13'b110000111000,
13'b110000111001,
13'b110001000001,
13'b110001000010,
13'b110001000011,
13'b110001000100,
13'b110001000101,
13'b110001000110,
13'b110001000111,
13'b110001001000,
13'b110001001001,
13'b110001001010,
13'b110001010001,
13'b110001010010,
13'b110001010011,
13'b110001010100,
13'b110001010101,
13'b110001010110,
13'b110001010111,
13'b110001011000,
13'b110001011001,
13'b110001011010,
13'b110001100001,
13'b110001100010,
13'b110001100011,
13'b110001100100,
13'b110001100101,
13'b110001100110,
13'b110001100111,
13'b110001101000,
13'b110001101001,
13'b110001101010,
13'b110001110001,
13'b110001110010,
13'b110001110011,
13'b110001110100,
13'b110001110101,
13'b110001110110,
13'b110001110111,
13'b110001111000,
13'b110001111001,
13'b110001111010,
13'b110010000001,
13'b110010000010,
13'b110010000011,
13'b110010000100,
13'b110010000101,
13'b110010000110,
13'b110010000111,
13'b110010001000,
13'b110010001001,
13'b110010001010,
13'b110010010010,
13'b110010010011,
13'b110010010100,
13'b110010010101,
13'b110010010110,
13'b110010010111,
13'b110010011010,
13'b110010100011,
13'b110010100100,
13'b110010100101,
13'b110010100110,
13'b110010100111,
13'b111000100011,
13'b111000100100,
13'b111000100101,
13'b111000110001,
13'b111000110010,
13'b111000110011,
13'b111000110100,
13'b111000110101,
13'b111000110110,
13'b111001000001,
13'b111001000010,
13'b111001000011,
13'b111001000100,
13'b111001000101,
13'b111001000110,
13'b111001000111,
13'b111001010001,
13'b111001010010,
13'b111001010011,
13'b111001010100,
13'b111001010101,
13'b111001010110,
13'b111001100001,
13'b111001100010,
13'b111001100011,
13'b111001100100,
13'b111001100101,
13'b111001100110,
13'b111001110001,
13'b111001110010,
13'b111001110011,
13'b111001110100,
13'b111001110101,
13'b111001110110,
13'b111010000010,
13'b111010000011,
13'b111010000100,
13'b111010000101,
13'b111010000110,
13'b111010010011,
13'b111010010100,
13'b111010010101,
13'b111010010110,
13'b111010100011,
13'b111010100100,
13'b111010100101,
13'b1000000110011,
13'b1000000110100,
13'b1000000110101,
13'b1000001000010,
13'b1000001000011,
13'b1000001000100,
13'b1000001000101,
13'b1000001010010,
13'b1000001010011,
13'b1000001010100,
13'b1000001010101,
13'b1000001100011,
13'b1000001100100,
13'b1000001100101,
13'b1000001110011,
13'b1000001110100,
13'b1000001110101,
13'b1000010000011,
13'b1000010000100,
13'b1000010000101,
13'b1000010010100,
13'b1000010010101,
13'b1001000110011,
13'b1001000110100,
13'b1001001000011,
13'b1001001000100,
13'b1001001010011,
13'b1001001010100,
13'b1001001100011,
13'b1001001100100: edge_mask_reg_512p3[510] <= 1'b1;
 		default: edge_mask_reg_512p3[510] <= 1'b0;
 	endcase

    case({x,y,z})
		default: edge_mask_reg_512p3[511] <= 1'b0;
 	endcase

end
endmodule

